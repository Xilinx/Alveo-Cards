/*
Copyright (c) 2023, Advanced Micro Devices, Inc. All rights reserved.
SPDX-License-Identifier: MIT
*/

//------------------------------------------------------------------------------

//
//  These compile flags are used for different configurations
//


`define CONFIG_FRAMES_TO_SEND 25
// Files: 
//       Sim/gtfmac_vnc_tb.v
// Usage:
//       Sets the number of frames to generate in the simulation.
