/*
Copyright (c) 2023, Advanced Micro Devices, Inc. All rights reserved.
SPDX-License-Identifier: MIT
*/

//------------------------------------------------------------------------------


//------{
`timescale 1fs/1fs
`default_nettype none
(* DowngradeIPIdentifiedWarnings="yes" *)
module gtfwizard_0_gtf_channel # (
  parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0,
  parameter [0:0] ACJTAG_MODE = 1'b0,
  parameter [0:0] ACJTAG_RESET = 1'b0,
  parameter [15:0] ADAPT_CFG0 = 16'h9200,
  parameter [15:0] ADAPT_CFG1 = 16'h801C,
  parameter [15:0] ADAPT_CFG2 = 16'h0000,
  parameter [0:0] A_RXOSCALRESET = 1'b0,
  parameter [0:0] A_RXPROGDIVRESET = 1'b0,
  parameter [0:0] A_RXTERMINATION = 1'b1,
  parameter [4:0] A_TXDIFFCTRL = 5'b01100,
  parameter [0:0] A_TXPROGDIVRESET = 1'b0,
  parameter CBCC_DATA_SOURCE_SEL = "DECODED",
  parameter [0:0] CDR_SWAP_MODE_EN = 1'b0,
  parameter [0:0] CFOK_PWRSVE_EN = 1'b1,
  parameter [15:0] CH_HSPMUX = 16'h2424,
  parameter [15:0] CKCAL1_CFG_0 = 16'b1100000011000000,
  parameter [15:0] CKCAL1_CFG_1 = 16'b0101000011000000,
  parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000,
  parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000,
  parameter [15:0] CKCAL2_CFG_0 = 16'b1100000011000000,
  parameter [15:0] CKCAL2_CFG_1 = 16'b1000000011000000,
  parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000,
  parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000,
  parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000,
  parameter [15:0] CPLL_CFG0 = 16'h01FA,
  parameter [15:0] CPLL_CFG1 = 16'h24A9,
  parameter [15:0] CPLL_CFG2 = 16'h6807,
  parameter [15:0] CPLL_CFG3 = 16'h0000,
  parameter integer CPLL_FBDIV = 4,
  parameter integer CPLL_FBDIV_45 = 4,
  parameter [15:0] CPLL_INIT_CFG0 = 16'h001E,
  parameter [15:0] CPLL_LOCK_CFG = 16'h01E8,
  parameter integer CPLL_REFCLK_DIV = 1,
  parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000,
  parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0,
  parameter [1:0] DDI_CTRL = 2'b00,
  parameter integer DDI_REALIGN_WAIT = 15,
  parameter [0:0] DELAY_ELEC = 1'b0,
  parameter [9:0] DMONITOR_CFG0 = 10'h000,
  parameter [7:0] DMONITOR_CFG1 = 8'h00,
  parameter [0:0] ES_CLK_PHASE_SEL = 1'b0,
  parameter [5:0] ES_CONTROL = 6'b000000,
  parameter ES_ERRDET_EN = "FALSE",
  parameter ES_EYE_SCAN_EN = "FALSE",
  parameter [11:0] ES_HORZ_OFFSET = 12'h800,
  parameter [4:0] ES_PRESCALE = 5'b00000,
  parameter [15:0] ES_QUALIFIER0 = 16'h0000,
  parameter [15:0] ES_QUALIFIER1 = 16'h0000,
  parameter [15:0] ES_QUALIFIER2 = 16'h0000,
  parameter [15:0] ES_QUALIFIER3 = 16'h0000,
  parameter [15:0] ES_QUALIFIER4 = 16'h0000,
  parameter [15:0] ES_QUALIFIER5 = 16'h0000,
  parameter [15:0] ES_QUALIFIER6 = 16'h0000,
  parameter [15:0] ES_QUALIFIER7 = 16'h0000,
  parameter [15:0] ES_QUALIFIER8 = 16'h0000,
  parameter [15:0] ES_QUALIFIER9 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK0 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK1 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK2 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK3 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK4 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK5 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK6 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK7 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK8 = 16'h0000,
  parameter [15:0] ES_QUAL_MASK9 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK0 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK1 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK2 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK3 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK4 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK5 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK6 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK7 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK8 = 16'h0000,
  parameter [15:0] ES_SDATA_MASK9 = 16'h0000,
  parameter integer EYESCAN_VP_RANGE = 0,
  parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0,
  parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111,
  parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111,
  parameter FTS_LANE_DESKEW_EN = "FALSE",
  parameter [4:0] GEARBOX_MODE = 5'b00000,
  parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0,
  parameter [0:0] LOCAL_MASTER = 1'b0,
  parameter integer LPBK_BIAS_CTRL = 4,
  parameter [0:0] LPBK_EN_RCAL_B = 1'b0,
  parameter [3:0] LPBK_EXT_RCAL = 4'b0000,
  parameter integer LPBK_IND_CTRL0 = 5,
  parameter integer LPBK_IND_CTRL1 = 5,
  parameter integer LPBK_IND_CTRL2 = 5,
  parameter integer LPBK_RG_CTRL = 2,
  parameter [15:0] MAC_CFG0 = 16'h0000,
  parameter [15:0] MAC_CFG1 = 16'h0000,
  parameter [15:0] MAC_CFG10 = 16'h00BB,
  parameter [15:0] MAC_CFG11 = 16'h0040,
  parameter [15:0] MAC_CFG12 = 16'h2580,
  parameter [15:0] MAC_CFG13 = 16'h0001,
  parameter [15:0] MAC_CFG14 = 16'h0000,
  parameter [15:0] MAC_CFG15 = 16'h0000,
  parameter [15:0] MAC_CFG2 = 16'h0000,
  parameter [15:0] MAC_CFG3 = 16'h0000,
  parameter [15:0] MAC_CFG4 = 16'h0000,
  parameter [15:0] MAC_CFG5 = 16'h0000,
  parameter [15:0] MAC_CFG6 = 16'h0000,
  parameter [15:0] MAC_CFG7 = 16'h0000,
  parameter [15:0] MAC_CFG8 = 16'h0000,
  parameter [15:0] MAC_CFG9 = 16'h0C03,
  parameter [15:0] PCS_RSVD0 = 16'h0000,
  parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C,
  parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19,
  parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64,
  parameter integer PREIQ_FREQ_BST = 0,
  parameter [15:0] RAW_MAC_CFG = 16'h0000,
  parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0,
  parameter [0:0] RCLK_SIPO_INV_EN = 1'b0,
  parameter [15:0] RCO_NEW_MAC_CFG0 = 16'h0000,
  parameter [15:0] RCO_NEW_MAC_CFG1 = 16'h0000,
  parameter [15:0] RCO_NEW_MAC_CFG2 = 16'h0000,
  parameter [15:0] RCO_NEW_MAC_CFG3 = 16'h0000,
  parameter [15:0] RCO_NEW_RAW_CFG0 = 16'h0000,
  parameter [15:0] RCO_NEW_RAW_CFG1 = 16'h2020,
  parameter [15:0] RCO_NEW_RAW_CFG2 = 16'h0000,
  parameter [15:0] RCO_NEW_RAW_CFG3 = 16'h0000,
  parameter [2:0] RTX_BUF_CML_CTRL = 3'b010,
  parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00,
  parameter [4:0] RXBUFRESET_TIME = 5'b00001,
  parameter RXBUF_EN = "TRUE",
  parameter [4:0] RXCDRFREQRESET_TIME = 5'b10000,
  parameter [4:0] RXCDRPHRESET_TIME = 5'b00001,
  parameter [15:0] RXCDR_CFG0 = 16'h0003,
  parameter [15:0] RXCDR_CFG1 = 16'h0000,
  parameter [15:0] RXCDR_CFG2 = 16'h0164,
  parameter [15:0] RXCDR_CFG3 = 16'h0024,
  parameter [15:0] RXCDR_CFG4 = 16'h5CF6,
  parameter [15:0] RXCDR_CFG5 = 16'hB46B,
  parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0,
  parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0,
  parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040,
  parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000,
  parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000,
  parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000,
  parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000,
  parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0,
  parameter [15:0] RXCFOK_CFG0 = 16'h0000,
  parameter [15:0] RXCFOK_CFG1 = 16'h0002,
  parameter [15:0] RXCFOK_CFG2 = 16'h002D,
  parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000,
  parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000,
  parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111,
  parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000,
  parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022,
  parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100,
  parameter [15:0] RXDFE_CFG0 = 16'h4000,
  parameter [15:0] RXDFE_CFG1 = 16'h0000,
  parameter [15:0] RXDFE_GC_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_GC_CFG1 = 16'h0000,
  parameter [15:0] RXDFE_GC_CFG2 = 16'h0000,
  parameter [15:0] RXDFE_H2_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H2_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H3_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H3_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H4_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H4_CFG1 = 16'h0003,
  parameter [15:0] RXDFE_H5_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H5_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H6_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H6_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H7_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H7_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H8_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H8_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_H9_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_H9_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HA_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HA_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HB_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HB_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HC_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HC_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HD_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HD_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HE_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HE_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_HF_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_HF_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_KH_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_KH_CFG1 = 16'h0000,
  parameter [15:0] RXDFE_KH_CFG2 = 16'h0000,
  parameter [15:0] RXDFE_KH_CFG3 = 16'h2000,
  parameter [15:0] RXDFE_OS_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_OS_CFG1 = 16'h0000,
  parameter [15:0] RXDFE_UT_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_UT_CFG1 = 16'h0002,
  parameter [15:0] RXDFE_UT_CFG2 = 16'h0000,
  parameter [15:0] RXDFE_VP_CFG0 = 16'h0000,
  parameter [15:0] RXDFE_VP_CFG1 = 16'h0022,
  parameter [15:0] RXDLY_CFG = 16'h0010,
  parameter [15:0] RXDLY_LCFG = 16'h0030,
  parameter [15:0] RXDLY_RAW_CFG = 16'h0010,
  parameter [15:0] RXDLY_RAW_LCFG = 16'h0000,
  parameter RXELECIDLE_CFG = "SIGCFG_4",
  parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4,
  parameter RXGEARBOX_EN = "FALSE",
  parameter [4:0] RXISCANRESET_TIME = 5'b00001,
  parameter [15:0] RXLPM_CFG = 16'h0000,
  parameter [15:0] RXLPM_GC_CFG = 16'h1000,
  parameter [15:0] RXLPM_KH_CFG0 = 16'h0000,
  parameter [15:0] RXLPM_KH_CFG1 = 16'h0002,
  parameter [15:0] RXLPM_OS_CFG0 = 16'h0000,
  parameter [15:0] RXLPM_OS_CFG1 = 16'h0000,
  parameter [4:0] RXOSCALRESET_TIME = 5'b00011,
  parameter integer RXOUT_DIV = 4,
  parameter [4:0] RXPCSRESET_TIME = 5'b00001,
  parameter [15:0] RXPHBEACON_CFG = 16'h0000,
  parameter [15:0] RXPHBEACON_RAW_CFG = 16'h0000,
  parameter [15:0] RXPHDLY_CFG = 16'h2020,
  parameter [15:0] RXPHSAMP_CFG = 16'h2100,
  parameter [15:0] RXPHSAMP_RAW_CFG = 16'h2100,
  parameter [15:0] RXPHSLIP_CFG = 16'h9933,
  parameter [15:0] RXPHSLIP_RAW_CFG = 16'h9933,
  parameter [4:0] RXPH_MONITOR_SEL = 5'b00000,
  parameter [15:0] RXPI_CFG0 = 16'h0102,
  parameter [15:0] RXPI_CFG1 = 16'b0000000001010100,
  parameter RXPMACLK_SEL = "DATA",
  parameter [4:0] RXPMARESET_TIME = 5'b00001,
  parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0,
  parameter integer RXPRBS_LINKACQ_CNT = 15,
  parameter [0:0] RXREFCLKDIV2_SEL = 1'b0,
  parameter integer RXSLIDE_AUTO_WAIT = 7,
  parameter RXSLIDE_MODE = "OFF",
  parameter [0:0] RXSYNC_MULTILANE = 1'b0,
  parameter [0:0] RXSYNC_OVRD = 1'b0,
  parameter [0:0] RXSYNC_SKIP_DA = 1'b0,
  parameter [0:0] RX_AFE_CM_EN = 1'b0,
  parameter [15:0] RX_BIAS_CFG0 = 16'h12B0,
  parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0,
  parameter integer RX_CLK25_DIV = 8,
  parameter [0:0] RX_CLKMUX_EN = 1'b1,
  parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000,
  parameter [3:0] RX_CM_BUF_CFG = 4'b1010,
  parameter [0:0] RX_CM_BUF_PD = 1'b0,
  parameter integer RX_CM_SEL = 2,
  parameter integer RX_CM_TRIM = 12,
  parameter [0:0] RX_CTLE_PWR_SAVING = 1'b0,
  parameter [3:0] RX_CTLE_RES_CTRL = 4'b0000,
  parameter integer RX_DATA_WIDTH = 20,
  parameter [5:0] RX_DDI_SEL = 6'b000000,
  parameter [2:0] RX_DEGEN_CTRL = 3'b100,
  parameter integer RX_DFELPM_CFG0 = 10,
  parameter [0:0] RX_DFELPM_CFG1 = 1'b1,
  parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1,
  parameter integer RX_DFE_AGC_CFG1 = 4,
  parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1,
  parameter integer RX_DFE_KL_LPM_KH_CFG1 = 2,
  parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01,
  parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4,
  parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0,
  parameter RX_DISPERR_SEQ_MATCH = "TRUE",
  parameter [4:0] RX_DIVRESET_TIME = 5'b00001,
  parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0,
  parameter integer RX_EN_SUM_RCAL_B = 0,
  parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000,
  parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0,
  parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b10,
  parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0,
  parameter [0:0] RX_I2V_FILTER_EN = 1'b1,
  parameter integer RX_INT_DATAWIDTH = 1,
  parameter [0:0] RX_PMA_POWER_SAVE = 1'b0,
  parameter [15:0] RX_PMA_RSV0 = 16'h002F,
  parameter real RX_PROGDIV_CFG = 0.0,
  parameter [15:0] RX_PROGDIV_RATE = 16'h0001,
  parameter [3:0] RX_RESLOAD_CTRL = 4'b0000,
  parameter [0:0] RX_RESLOAD_OVRD = 1'b0,
  parameter [2:0] RX_SAMPLE_PERIOD = 3'b101,
  parameter integer RX_SIG_VALID_DLY = 11,
  parameter integer RX_SUM_DEGEN_AVTT_OVERITE = 0,
  parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0,
  parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000,
  parameter integer RX_SUM_PWR_SAVING = 0,
  parameter [3:0] RX_SUM_RES_CTRL = 4'b0000,
  parameter [3:0] RX_SUM_VCMTUNE = 4'b0011,
  parameter [0:0] RX_SUM_VCM_BIAS_TUNE_EN = 1'b1,
  parameter [0:0] RX_SUM_VCM_OVWR = 1'b0,
  parameter [2:0] RX_SUM_VREF_TUNE = 3'b100,
  parameter [1:0] RX_TUNE_AFE_OS = 2'b00,
  parameter [2:0] RX_VREG_CTRL = 3'b010,
  parameter [0:0] RX_VREG_PDB = 1'b1,
  parameter [1:0] RX_WIDEMODE_CDR = 2'b01,
  parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01,
  parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01,
  parameter RX_XCLK_SEL = "RXDES",
  parameter [0:0] RX_XMODE_SEL = 1'b0,
  parameter [0:0] SAMPLE_CLK_PHASE = 1'b0,
  parameter SATA_CPLL_CFG = "VCO_3000MHZ",
  parameter SIM_MODE = "FAST",
  parameter SIM_RESET_SPEEDUP = "TRUE",
  parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z",
  parameter [0:0] SRSTMODE = 1'b0,
  parameter [1:0] TAPDLY_SET_TX = 2'h0,
  parameter [15:0] TCO_NEW_CFG0 = 16'h0000,
  parameter [15:0] TCO_NEW_CFG1 = 16'h0000,
  parameter [15:0] TCO_NEW_CFG2 = 16'h0000,
  parameter [15:0] TCO_NEW_CFG3 = 16'h0000,
  parameter [15:0] TCO_RSVD1 = 16'h0000,
  parameter [15:0] TCO_RSVD2 = 16'h0000,
  parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000,
  parameter [2:0] TERM_RCAL_OVRD = 3'b000,
  parameter [7:0] TRANS_TIME_RATE = 8'h0E,
  parameter [7:0] TST_RSV0 = 8'h00,
  parameter [7:0] TST_RSV1 = 8'h00,
  parameter TXBUF_EN = "TRUE",
  parameter [15:0] TXDLY_CFG = 16'h0010,
  parameter [15:0] TXDLY_LCFG = 16'h0030,
  parameter integer TXDRV_FREQBAND = 0,
  parameter [15:0] TXFE_CFG0 = 16'h0000,
  parameter [15:0] TXFE_CFG1 = 16'h0000,
  parameter [15:0] TXFE_CFG2 = 16'h0000,
  parameter [15:0] TXFE_CFG3 = 16'h0000,
  parameter TXFIFO_ADDR_CFG = "LOW",
  parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4,
  parameter integer TXOUT_DIV = 4,
  parameter [4:0] TXPCSRESET_TIME = 5'b00001,
  parameter [15:0] TXPHDLY_CFG0 = 16'h6020,
  parameter [15:0] TXPHDLY_CFG1 = 16'h0002,
  parameter [15:0] TXPH_CFG = 16'h0103,
  parameter [15:0] TXPH_CFG2 = 16'h0000,
  parameter [4:0] TXPH_MONITOR_SEL = 5'b00000,
  parameter [15:0] TXPI_CFG0 = 16'h0100,
  parameter [15:0] TXPI_CFG1 = 16'h0000,
  parameter [0:0] TXPI_GRAY_SEL = 1'b0,
  parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0,
  parameter [0:0] TXPI_PPM = 1'b0,
  parameter [7:0] TXPI_PPM_CFG = 8'b00000000,
  parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000,
  parameter [4:0] TXPMARESET_TIME = 5'b00001,
  parameter [0:0] TXREFCLKDIV2_SEL = 1'b0,
  parameter integer TXSWBST_BST = 1,
  parameter integer TXSWBST_EN = 0,
  parameter integer TXSWBST_MAG = 6,
  parameter [0:0] TXSYNC_MULTILANE = 1'b0,
  parameter [0:0] TXSYNC_OVRD = 1'b0,
  parameter [0:0] TXSYNC_SKIP_DA = 1'b0,
  parameter integer TX_CLK25_DIV = 8,
  parameter [0:0] TX_CLKMUX_EN = 1'b1,
  parameter integer TX_DATA_WIDTH = 20,
  parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000,
  parameter [4:0] TX_DIVRESET_TIME = 5'b00001,
  parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110,
  parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100,
  parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0,
  parameter [0:0] TX_FIFO_BYP_EN = 1'b0,
  parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0,
  parameter integer TX_INT_DATAWIDTH = 0,
  parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE",
  parameter [0:0] TX_MAINCURSOR_SEL = 1'b0,
  parameter [15:0] TX_PHICAL_CFG0 = 16'h0000,
  parameter [15:0] TX_PHICAL_CFG1 = 16'h003F,
  parameter integer TX_PI_BIASSET = 0,
  parameter [0:0] TX_PMADATA_OPT = 1'b0,
  parameter [0:0] TX_PMA_POWER_SAVE = 1'b0,
  parameter [15:0] TX_PMA_RSV0 = 16'h0000,
  parameter [15:0] TX_PMA_RSV1 = 16'h0000,
  parameter TX_PROGCLK_SEL = "POSTPI",
  parameter real TX_PROGDIV_CFG = 0.0,
  parameter [15:0] TX_PROGDIV_RATE = 16'h0001,
  parameter [2:0] TX_SAMPLE_PERIOD = 3'b101,
  parameter [1:0] TX_SW_MEAS = 2'b00,
  parameter [2:0] TX_VREG_CTRL = 3'b000,
  parameter [0:0] TX_VREG_PDB = 1'b0,
  parameter [1:0] TX_VREG_VREFSEL = 2'b00,
  parameter TX_XCLK_SEL = "TXOUT",
  parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0,
  parameter [0:0] USE_RAW_ELEC = 1'b0,
  parameter [0:0] Y_ALL_MODE = 1'b0
)(
  input  wire   gtf_ch_cdrstepdir,
  input  wire   gtf_ch_cdrstepsq,
  input  wire   gtf_ch_cdrstepsx,
  input  wire   gtf_ch_cfgreset,
  input  wire   gtf_ch_clkrsvd0,
  input  wire   gtf_ch_clkrsvd1,
  input  wire   gtf_ch_cpllfreqlock,
  input  wire   gtf_ch_cplllockdetclk,
  input  wire   gtf_ch_cplllocken,
  input  wire   gtf_ch_cpllpd,
  input  wire   gtf_ch_cpllreset,
  input  wire   gtf_ch_ctltxresendpause,
  input  wire   gtf_ch_ctltxsendidle,
  input  wire   gtf_ch_ctltxsendlfi,
  input  wire   gtf_ch_ctltxsendrfi,
  input  wire   gtf_ch_dmonfiforeset,
  input  wire   gtf_ch_dmonitorclk,
  input  wire   gtf_ch_drpclk,
  input  wire   gtf_ch_drpen,
  input  wire   gtf_ch_drprst,
  input  wire   gtf_ch_drpwe,
  input  wire   gtf_ch_eyescanreset,
  input  wire   gtf_ch_eyescantrigger,
  input  wire   gtf_ch_freqos,
  input  wire   gtf_ch_gtfrxn,
  input  wire   gtf_ch_gtfrxp,
  input  wire   gtf_ch_gtgrefclk,
  input  wire   gtf_ch_gtnorthrefclk0,
  input  wire   gtf_ch_gtnorthrefclk1,
  input  wire   gtf_ch_gtrefclk0,
  input  wire   gtf_ch_gtrefclk1,
  input  wire   gtf_ch_gtrxreset,
  input  wire   gtf_ch_gtrxresetsel,
  input  wire   gtf_ch_gtsouthrefclk0,
  input  wire   gtf_ch_gtsouthrefclk1,
  input  wire   gtf_ch_gttxreset,
  input  wire   gtf_ch_gttxresetsel,
  input  wire   gtf_ch_incpctrl,
  input  wire   gtf_ch_qpll0clk,
  input  wire   gtf_ch_qpll0freqlock,
  input  wire   gtf_ch_qpll0refclk,
  input  wire   gtf_ch_qpll1clk,
  input  wire   gtf_ch_qpll1freqlock,
  input  wire   gtf_ch_qpll1refclk,
  input  wire   gtf_ch_resetovrd,
  input  wire   gtf_ch_rxafecfoken,
  input  wire   gtf_ch_rxcdrfreqreset,
  input  wire   gtf_ch_rxcdrhold,
  input  wire   gtf_ch_rxcdrovrden,
  input  wire   gtf_ch_rxcdrreset,
  input  wire   gtf_ch_rxckcalreset,
  input  wire   gtf_ch_rxdfeagchold,
  input  wire   gtf_ch_rxdfeagcovrden,
  input  wire   gtf_ch_rxdfecfokfen,
  input  wire   gtf_ch_rxdfecfokfpulse,
  input  wire   gtf_ch_rxdfecfokhold,
  input  wire   gtf_ch_rxdfecfokovren,
  input  wire   gtf_ch_rxdfekhhold,
  input  wire   gtf_ch_rxdfekhovrden,
  input  wire   gtf_ch_rxdfelfhold,
  input  wire   gtf_ch_rxdfelfovrden,
  input  wire   gtf_ch_rxdfelpmreset,
  input  wire   gtf_ch_rxdfetap10hold,
  input  wire   gtf_ch_rxdfetap10ovrden,
  input  wire   gtf_ch_rxdfetap11hold,
  input  wire   gtf_ch_rxdfetap11ovrden,
  input  wire   gtf_ch_rxdfetap12hold,
  input  wire   gtf_ch_rxdfetap12ovrden,
  input  wire   gtf_ch_rxdfetap13hold,
  input  wire   gtf_ch_rxdfetap13ovrden,
  input  wire   gtf_ch_rxdfetap14hold,
  input  wire   gtf_ch_rxdfetap14ovrden,
  input  wire   gtf_ch_rxdfetap15hold,
  input  wire   gtf_ch_rxdfetap15ovrden,
  input  wire   gtf_ch_rxdfetap2hold,
  input  wire   gtf_ch_rxdfetap2ovrden,
  input  wire   gtf_ch_rxdfetap3hold,
  input  wire   gtf_ch_rxdfetap3ovrden,
  input  wire   gtf_ch_rxdfetap4hold,
  input  wire   gtf_ch_rxdfetap4ovrden,
  input  wire   gtf_ch_rxdfetap5hold,
  input  wire   gtf_ch_rxdfetap5ovrden,
  input  wire   gtf_ch_rxdfetap6hold,
  input  wire   gtf_ch_rxdfetap6ovrden,
  input  wire   gtf_ch_rxdfetap7hold,
  input  wire   gtf_ch_rxdfetap7ovrden,
  input  wire   gtf_ch_rxdfetap8hold,
  input  wire   gtf_ch_rxdfetap8ovrden,
  input  wire   gtf_ch_rxdfetap9hold,
  input  wire   gtf_ch_rxdfetap9ovrden,
  input  wire   gtf_ch_rxdfeuthold,
  input  wire   gtf_ch_rxdfeutovrden,
  input  wire   gtf_ch_rxdfevphold,
  input  wire   gtf_ch_rxdfevpovrden,
  input  wire   gtf_ch_rxdfexyden,
  input  wire   gtf_ch_rxdlybypass,
  input  wire   gtf_ch_rxdlyen,
  input  wire   gtf_ch_rxdlyovrden,
  input  wire   gtf_ch_rxdlysreset,
  input  wire   gtf_ch_rxlpmen,
  input  wire   gtf_ch_rxlpmgchold,
  input  wire   gtf_ch_rxlpmgcovrden,
  input  wire   gtf_ch_rxlpmhfhold,
  input  wire   gtf_ch_rxlpmhfovrden,
  input  wire   gtf_ch_rxlpmlfhold,
  input  wire   gtf_ch_rxlpmlfklovrden,
  input  wire   gtf_ch_rxlpmoshold,
  input  wire   gtf_ch_rxlpmosovrden,
  input  wire   gtf_ch_rxoscalreset,
  input  wire   gtf_ch_rxoshold,
  input  wire   gtf_ch_rxosovrden,
  input  wire   gtf_ch_rxpcsreset,
  input  wire   gtf_ch_rxphalign,
  input  wire   gtf_ch_rxphalignen,
  input  wire   gtf_ch_rxphdlypd,
  input  wire   gtf_ch_rxphdlyreset,
  input  wire   gtf_ch_rxpmareset,
  input  wire   gtf_ch_rxpolarity,
  input  wire   gtf_ch_rxprbscntreset,
  input  wire   gtf_ch_rxprogdivreset,
  input  wire   gtf_ch_rxslipoutclk,
  input  wire   gtf_ch_rxslippma,
  input  wire   gtf_ch_rxsyncallin,
  input  wire   gtf_ch_rxsyncin,
  input  wire   gtf_ch_rxsyncmode,
  input  wire   gtf_ch_rxtermination,
  input  wire   gtf_ch_rxuserrdy,
  input  wire   gtf_ch_rxusrclk,
  input  wire   gtf_ch_rxusrclk2,
  input  wire   gtf_ch_txaxisterr,
  input  wire   gtf_ch_txaxistpoison,
  input  wire   gtf_ch_txaxistvalid,
  input  wire   gtf_ch_txdccforcestart,
  input  wire   gtf_ch_txdccreset,
  input  wire   gtf_ch_txdlybypass,
  input  wire   gtf_ch_txdlyen,
  input  wire   gtf_ch_txdlyhold,
  input  wire   gtf_ch_txdlyovrden,
  input  wire   gtf_ch_txdlysreset,
  input  wire   gtf_ch_txdlyupdown,
  input  wire   gtf_ch_txelecidle,
  input  wire   gtf_ch_txgbseqsync,
  input  wire   gtf_ch_txmuxdcdexhold,
  input  wire   gtf_ch_txmuxdcdorwren,
  input  wire   gtf_ch_txpcsreset,
  input  wire   gtf_ch_txphalign,
  input  wire   gtf_ch_txphalignen,
  input  wire   gtf_ch_txphdlypd,
  input  wire   gtf_ch_txphdlyreset,
  input  wire   gtf_ch_txphdlytstclk,
  input  wire   gtf_ch_txphinit,
  input  wire   gtf_ch_txphovrden,
  input  wire   gtf_ch_txpippmen,
  input  wire   gtf_ch_txpippmovrden,
  input  wire   gtf_ch_txpippmpd,
  input  wire   gtf_ch_txpippmsel,
  input  wire   gtf_ch_txpisopd,
  input  wire   gtf_ch_txpmareset,
  input  wire   gtf_ch_txpolarity,
  input  wire   gtf_ch_txprbsforceerr,
  input  wire   gtf_ch_txprogdivreset,
  input  wire   gtf_ch_txsyncallin,
  input  wire   gtf_ch_txsyncin,
  input  wire   gtf_ch_txsyncmode,
  input  wire   gtf_ch_txuserrdy,
  input  wire   gtf_ch_txusrclk,
  input  wire   gtf_ch_txusrclk2,
  input  wire [15:0]  gtf_ch_drpdi,
  input  wire [15:0]  gtf_ch_gtrsvd,
  input  wire [15:0]  gtf_ch_pcsrsvdin,
  input  wire [19:0]  gtf_ch_tstin,
  input  wire [1:0]   gtf_ch_rxelecidlemode,
  input  wire [1:0]   gtf_ch_rxmonitorsel,
  input  wire [1:0]   gtf_ch_rxpd,
  input  wire [1:0]   gtf_ch_rxpllclksel,
  input  wire [1:0]   gtf_ch_rxsysclksel,
  input  wire [1:0]   gtf_ch_txaxistsof,
  input  wire [1:0]   gtf_ch_txpd,
  input  wire [1:0]   gtf_ch_txpllclksel,
  input  wire [1:0]   gtf_ch_txsysclksel,
  input  wire [2:0]   gtf_ch_cpllrefclksel,
  input  wire [2:0]   gtf_ch_loopback,
  input  wire [2:0]   gtf_ch_rxoutclksel,
  input  wire [2:0]   gtf_ch_txoutclksel,
  input  wire [39:0]  gtf_ch_txrawdata,
  input  wire [3:0]   gtf_ch_rxdfecfokfcnum,
  input  wire [3:0]   gtf_ch_rxprbssel,
  input  wire [3:0]   gtf_ch_txprbssel,
  input  wire [4:0]   gtf_ch_txaxistterm,
  input  wire [4:0]   gtf_ch_txdiffctrl,
  input  wire [4:0]   gtf_ch_txpippmstepsize,
  input  wire [4:0]   gtf_ch_txpostcursor,
  input  wire [4:0]   gtf_ch_txprecursor,
  input  wire [63:0]  gtf_ch_txaxistdata,
  input  wire [6:0]   gtf_ch_rxckcalstart,
  input  wire [6:0]   gtf_ch_txmaincursor,
  input  wire [7:0]   gtf_ch_txaxistlast,
  input  wire [7:0]   gtf_ch_txaxistpre,
  input  wire [8:0]   gtf_ch_ctlrxpauseack,
  input  wire [8:0]   gtf_ch_ctltxpausereq,
  input  wire [9:0]   gtf_ch_drpaddr,
  output wire       gtf_ch_cpllfbclklost,
  output wire       gtf_ch_cplllock,
  output wire       gtf_ch_cpllrefclklost,
  output wire       gtf_ch_dmonitoroutclk,
  output wire       gtf_ch_drprdy,
  output wire       gtf_ch_eyescandataerror,
  output wire       gtf_ch_gtftxn,
  output wire       gtf_ch_gtftxp,
  output wire       gtf_ch_gtpowergood,
  output wire       gtf_ch_gtrefclkmonitor,
  output wire       gtf_ch_resetexception,
  output wire       gtf_ch_rxaxisterr,
  output wire       gtf_ch_rxaxistvalid,
  output wire       gtf_ch_rxbitslip,
  output wire       gtf_ch_rxcdrlock,
  output wire       gtf_ch_rxcdrphdone,
  output wire       gtf_ch_rxckcaldone,
  output wire       gtf_ch_rxdlysresetdone,
  output wire       gtf_ch_rxelecidle,
  output wire       gtf_ch_rxgbseqstart,
  output wire       gtf_ch_rxosintdone,
  output wire       gtf_ch_rxosintstarted,
  output wire       gtf_ch_rxosintstrobedone,
  output wire       gtf_ch_rxosintstrobestarted,
  output wire       gtf_ch_rxoutclk,
  output wire       gtf_ch_rxoutclkfabric,
  output wire       gtf_ch_rxoutclkpcs,
  output wire       gtf_ch_rxphaligndone,
  output wire       gtf_ch_rxphalignerr,
  output wire       gtf_ch_rxpmaresetdone,
  output wire       gtf_ch_rxprbserr,
  output wire       gtf_ch_rxprbslocked,
  output wire       gtf_ch_rxprgdivresetdone,
  output wire       gtf_ch_rxptpsop,
  output wire       gtf_ch_rxptpsoppos,
  output wire       gtf_ch_rxrecclkout,
  output wire       gtf_ch_rxresetdone,
  output wire       gtf_ch_rxslipdone,
  output wire       gtf_ch_rxslipoutclkrdy,
  output wire       gtf_ch_rxslippmardy,
  output wire       gtf_ch_rxsyncdone,
  output wire       gtf_ch_rxsyncout,
  output wire       gtf_ch_statrxbadcode,
  output wire       gtf_ch_statrxbadfcs,
  output wire       gtf_ch_statrxbadpreamble,
  output wire       gtf_ch_statrxbadsfd,
  output wire       gtf_ch_statrxblocklock,
  output wire       gtf_ch_statrxbroadcast,
  output wire       gtf_ch_statrxfcserr,
  output wire       gtf_ch_statrxframingerr,
  output wire       gtf_ch_statrxgotsignalos,
  output wire       gtf_ch_statrxhiber,
  output wire       gtf_ch_statrxinrangeerr,
  output wire       gtf_ch_statrxinternallocalfault,
  output wire       gtf_ch_statrxlocalfault,
  output wire       gtf_ch_statrxmulticast,
  output wire       gtf_ch_statrxpkt,
  output wire       gtf_ch_statrxpkterr,
  output wire       gtf_ch_statrxreceivedlocalfault,
  output wire       gtf_ch_statrxremotefault,
  output wire       gtf_ch_statrxstatus,
  output wire       gtf_ch_statrxstompedfcs,
  output wire       gtf_ch_statrxtestpatternmismatch,
  output wire       gtf_ch_statrxtruncated,
  output wire       gtf_ch_statrxunicast,
  output wire       gtf_ch_statrxvalidctrlcode,
  output wire       gtf_ch_statrxvlan,
  output wire       gtf_ch_stattxbadfcs,
  output wire       gtf_ch_stattxbroadcast,
  output wire       gtf_ch_stattxfcserr,
  output wire       gtf_ch_stattxmulticast,
  output wire       gtf_ch_stattxpkt,
  output wire       gtf_ch_stattxpkterr,
  output wire       gtf_ch_stattxunicast,
  output wire       gtf_ch_stattxvlan,
  output wire       gtf_ch_txaxistready,
  output wire       gtf_ch_txdccdone,
  output wire       gtf_ch_txdlysresetdone,
  output wire       gtf_ch_txgbseqstart,
  output wire       gtf_ch_txoutclk,
  output wire       gtf_ch_txoutclkfabric,
  output wire       gtf_ch_txoutclkpcs,
  output wire       gtf_ch_txphaligndone,
  output wire       gtf_ch_txphinitdone,
  output wire       gtf_ch_txpmaresetdone,
  output wire       gtf_ch_txprgdivresetdone,
  output wire       gtf_ch_txptpsop,
  output wire       gtf_ch_txptpsoppos,
  output wire       gtf_ch_txresetdone,
  output wire       gtf_ch_txsyncdone,
  output wire       gtf_ch_txsyncout,
  output wire       gtf_ch_txunfout,
  output wire [15:0] gtf_ch_dmonitorout,
  output wire [15:0] gtf_ch_drpdo,
  output wire [15:0] gtf_ch_pcsrsvdout,
  output wire [15:0] gtf_ch_pinrsrvdas,
  output wire [1:0]  gtf_ch_rxaxistsof,
  output wire [39:0] gtf_ch_rxrawdata,
  output wire [3:0]  gtf_ch_statrxbytes,
  output wire [3:0]  gtf_ch_stattxbytes,
  output wire [4:0]  gtf_ch_rxaxistterm,
  output wire [63:0] gtf_ch_rxaxistdata,
  output wire [7:0]  gtf_ch_rxaxistlast,
  output wire [7:0]  gtf_ch_rxaxistpre,
  output wire [7:0]  gtf_ch_rxmonitorout,
  output wire [8:0]  gtf_ch_statrxpausequanta,
  output wire [8:0]  gtf_ch_statrxpausereq,
  output wire [8:0]  gtf_ch_statrxpausevalid,
  output wire [8:0]  gtf_ch_stattxpausevalid
);


//----{
GTF_CHANNEL #(
.ACJTAG_DEBUG_MODE             (ACJTAG_DEBUG_MODE              ),
.ACJTAG_MODE                   (ACJTAG_MODE                    ),
.ACJTAG_RESET                  (ACJTAG_RESET                   ),
.ADAPT_CFG0                    (ADAPT_CFG0                     ),
.ADAPT_CFG1                    (ADAPT_CFG1                     ),
.ADAPT_CFG2                    (ADAPT_CFG2                     ),
.A_RXOSCALRESET                (A_RXOSCALRESET                 ),
.A_RXPROGDIVRESET              (A_RXPROGDIVRESET               ),
.A_RXTERMINATION               (A_RXTERMINATION                ),
.A_TXDIFFCTRL                  (A_TXDIFFCTRL                   ),
.A_TXPROGDIVRESET              (A_TXPROGDIVRESET               ),
.CBCC_DATA_SOURCE_SEL          (CBCC_DATA_SOURCE_SEL           ),
.CDR_SWAP_MODE_EN              (CDR_SWAP_MODE_EN               ),
.CFOK_PWRSVE_EN                (CFOK_PWRSVE_EN                 ),
.CH_HSPMUX                     (CH_HSPMUX                      ),
.CKCAL1_CFG_0                  (CKCAL1_CFG_0                   ),
.CKCAL1_CFG_1                  (CKCAL1_CFG_1                   ),
.CKCAL1_CFG_2                  (CKCAL1_CFG_2                   ),
.CKCAL1_CFG_3                  (CKCAL1_CFG_3                   ),
.CKCAL2_CFG_0                  (CKCAL2_CFG_0                   ),
.CKCAL2_CFG_1                  (CKCAL2_CFG_1                   ),
.CKCAL2_CFG_2                  (CKCAL2_CFG_2                   ),
.CKCAL2_CFG_3                  (CKCAL2_CFG_3                   ),
.CKCAL2_CFG_4                  (CKCAL2_CFG_4                   ),
.CPLL_CFG0                     (CPLL_CFG0                      ),
.CPLL_CFG1                     (CPLL_CFG1                      ),
.CPLL_CFG2                     (CPLL_CFG2                      ),
.CPLL_CFG3                     (CPLL_CFG3                      ),
.CPLL_FBDIV                    (CPLL_FBDIV                     ),
.CPLL_FBDIV_45                 (CPLL_FBDIV_45                  ),
.CPLL_INIT_CFG0                (CPLL_INIT_CFG0                 ),
.CPLL_LOCK_CFG                 (CPLL_LOCK_CFG                  ),
.CPLL_REFCLK_DIV               (CPLL_REFCLK_DIV                ),
.CTLE3_OCAP_EXT_CTRL           (CTLE3_OCAP_EXT_CTRL            ),
.CTLE3_OCAP_EXT_EN             (CTLE3_OCAP_EXT_EN              ),
.DDI_CTRL                      (DDI_CTRL                       ),
.DDI_REALIGN_WAIT              (DDI_REALIGN_WAIT               ),
.DELAY_ELEC                    (DELAY_ELEC                     ),
.DMONITOR_CFG0                 (DMONITOR_CFG0                  ),
.DMONITOR_CFG1                 (DMONITOR_CFG1                  ),
.ES_CLK_PHASE_SEL              (ES_CLK_PHASE_SEL               ),
.ES_CONTROL                    (ES_CONTROL                     ),
.ES_ERRDET_EN                  (ES_ERRDET_EN                   ),
.ES_EYE_SCAN_EN                (ES_EYE_SCAN_EN                 ),
.ES_HORZ_OFFSET                (ES_HORZ_OFFSET                 ),
.ES_PRESCALE                   (ES_PRESCALE                    ),
.ES_QUALIFIER0                 (ES_QUALIFIER0                  ),
.ES_QUALIFIER1                 (ES_QUALIFIER1                  ),
.ES_QUALIFIER2                 (ES_QUALIFIER2                  ),
.ES_QUALIFIER3                 (ES_QUALIFIER3                  ),
.ES_QUALIFIER4                 (ES_QUALIFIER4                  ),
.ES_QUALIFIER5                 (ES_QUALIFIER5                  ),
.ES_QUALIFIER6                 (ES_QUALIFIER6                  ),
.ES_QUALIFIER7                 (ES_QUALIFIER7                  ),
.ES_QUALIFIER8                 (ES_QUALIFIER8                  ),
.ES_QUALIFIER9                 (ES_QUALIFIER9                  ),
.ES_QUAL_MASK0                 (ES_QUAL_MASK0                  ),
.ES_QUAL_MASK1                 (ES_QUAL_MASK1                  ),
.ES_QUAL_MASK2                 (ES_QUAL_MASK2                  ),
.ES_QUAL_MASK3                 (ES_QUAL_MASK3                  ),
.ES_QUAL_MASK4                 (ES_QUAL_MASK4                  ),
.ES_QUAL_MASK5                 (ES_QUAL_MASK5                  ),
.ES_QUAL_MASK6                 (ES_QUAL_MASK6                  ),
.ES_QUAL_MASK7                 (ES_QUAL_MASK7                  ),
.ES_QUAL_MASK8                 (ES_QUAL_MASK8                  ),
.ES_QUAL_MASK9                 (ES_QUAL_MASK9                  ),
.ES_SDATA_MASK0                (ES_SDATA_MASK0                 ),
.ES_SDATA_MASK1                (ES_SDATA_MASK1                 ),
.ES_SDATA_MASK2                (ES_SDATA_MASK2                 ),
.ES_SDATA_MASK3                (ES_SDATA_MASK3                 ),
.ES_SDATA_MASK4                (ES_SDATA_MASK4                 ),
.ES_SDATA_MASK5                (ES_SDATA_MASK5                 ),
.ES_SDATA_MASK6                (ES_SDATA_MASK6                 ),
.ES_SDATA_MASK7                (ES_SDATA_MASK7                 ),
.ES_SDATA_MASK8                (ES_SDATA_MASK8                 ),
.ES_SDATA_MASK9                (ES_SDATA_MASK9                 ),
.EYESCAN_VP_RANGE              (EYESCAN_VP_RANGE               ),
.EYE_SCAN_SWAP_EN              (EYE_SCAN_SWAP_EN               ),
.FTS_DESKEW_SEQ_ENABLE         (FTS_DESKEW_SEQ_ENABLE          ),
.FTS_LANE_DESKEW_CFG           (FTS_LANE_DESKEW_CFG            ),
.FTS_LANE_DESKEW_EN            (FTS_LANE_DESKEW_EN             ),
.GEARBOX_MODE                  (GEARBOX_MODE                   ),
.ISCAN_CK_PH_SEL2              (ISCAN_CK_PH_SEL2               ),
.LOCAL_MASTER                  (LOCAL_MASTER                   ),
.LPBK_BIAS_CTRL                (LPBK_BIAS_CTRL                 ),
.LPBK_EN_RCAL_B                (LPBK_EN_RCAL_B                 ),
.LPBK_EXT_RCAL                 (LPBK_EXT_RCAL                  ),
.LPBK_IND_CTRL0                (LPBK_IND_CTRL0                 ),
.LPBK_IND_CTRL1                (LPBK_IND_CTRL1                 ),
.LPBK_IND_CTRL2                (LPBK_IND_CTRL2                 ),
.LPBK_RG_CTRL                  (LPBK_RG_CTRL                   ),
.MAC_CFG0                      (MAC_CFG0                       ),
.MAC_CFG1                      (MAC_CFG1                       ),
.MAC_CFG10                     (MAC_CFG10                      ),
.MAC_CFG11                     (MAC_CFG11                      ),
.MAC_CFG12                     (MAC_CFG12                      ),
.MAC_CFG13                     (MAC_CFG13                      ),
.MAC_CFG14                     (MAC_CFG14                      ),
.MAC_CFG15                     (MAC_CFG15                      ),
.MAC_CFG2                      (MAC_CFG2                       ),
.MAC_CFG3                      (MAC_CFG3                       ),
.MAC_CFG4                      (MAC_CFG4                       ),
.MAC_CFG5                      (MAC_CFG5                       ),
.MAC_CFG6                      (MAC_CFG6                       ),
.MAC_CFG7                      (MAC_CFG7                       ),
.MAC_CFG8                      (MAC_CFG8                       ),
.MAC_CFG9                      (MAC_CFG9                       ),
.PCS_RSVD0                     (PCS_RSVD0                      ),
.PD_TRANS_TIME_FROM_P2         (PD_TRANS_TIME_FROM_P2          ),
.PD_TRANS_TIME_NONE_P2         (PD_TRANS_TIME_NONE_P2          ),
.PD_TRANS_TIME_TO_P2           (PD_TRANS_TIME_TO_P2            ),
.PREIQ_FREQ_BST                (PREIQ_FREQ_BST                 ),
.RAW_MAC_CFG                   (RAW_MAC_CFG                    ),
.RCLK_SIPO_DLY_ENB             (RCLK_SIPO_DLY_ENB              ),
.RCLK_SIPO_INV_EN              (RCLK_SIPO_INV_EN               ),
.RCO_NEW_MAC_CFG0              (RCO_NEW_MAC_CFG0               ),
.RCO_NEW_MAC_CFG1              (RCO_NEW_MAC_CFG1               ),
.RCO_NEW_MAC_CFG2              (RCO_NEW_MAC_CFG2               ),
.RCO_NEW_MAC_CFG3              (RCO_NEW_MAC_CFG3               ),
.RCO_NEW_RAW_CFG0              (RCO_NEW_RAW_CFG0               ),
.RCO_NEW_RAW_CFG1              (RCO_NEW_RAW_CFG1               ),
.RCO_NEW_RAW_CFG2              (RCO_NEW_RAW_CFG2               ),
.RCO_NEW_RAW_CFG3              (RCO_NEW_RAW_CFG3               ),
.RTX_BUF_CML_CTRL              (RTX_BUF_CML_CTRL               ),
.RTX_BUF_TERM_CTRL             (RTX_BUF_TERM_CTRL              ),
.RXBUFRESET_TIME               (RXBUFRESET_TIME                ),
.RXBUF_EN                      (RXBUF_EN                       ),
.RXCDRFREQRESET_TIME           (RXCDRFREQRESET_TIME            ),
.RXCDRPHRESET_TIME             (RXCDRPHRESET_TIME              ),
.RXCDR_CFG0                    (RXCDR_CFG0                     ),
.RXCDR_CFG1                    (RXCDR_CFG1                     ),
.RXCDR_CFG2                    (RXCDR_CFG2                     ),
.RXCDR_CFG3                    (RXCDR_CFG3                     ),
.RXCDR_CFG4                    (RXCDR_CFG4                     ),
.RXCDR_CFG5                    (RXCDR_CFG5                     ),
.RXCDR_FR_RESET_ON_EIDLE       (RXCDR_FR_RESET_ON_EIDLE        ),
.RXCDR_HOLD_DURING_EIDLE       (RXCDR_HOLD_DURING_EIDLE        ),
.RXCDR_LOCK_CFG0               (RXCDR_LOCK_CFG0                ),
.RXCDR_LOCK_CFG1               (RXCDR_LOCK_CFG1                ),
.RXCDR_LOCK_CFG2               (RXCDR_LOCK_CFG2                ),
.RXCDR_LOCK_CFG3               (RXCDR_LOCK_CFG3                ),
.RXCDR_LOCK_CFG4               (RXCDR_LOCK_CFG4                ),
.RXCDR_PH_RESET_ON_EIDLE       (RXCDR_PH_RESET_ON_EIDLE        ),
.RXCFOK_CFG0                   (RXCFOK_CFG0                    ),
.RXCFOK_CFG1                   (RXCFOK_CFG1                    ),
.RXCFOK_CFG2                   (RXCFOK_CFG2                    ),
.RXCKCAL1_IQ_LOOP_RST_CFG      (RXCKCAL1_IQ_LOOP_RST_CFG       ),
.RXCKCAL1_I_LOOP_RST_CFG       (RXCKCAL1_I_LOOP_RST_CFG        ),
.RXCKCAL1_Q_LOOP_RST_CFG       (RXCKCAL1_Q_LOOP_RST_CFG        ),
.RXCKCAL2_DX_LOOP_RST_CFG      (RXCKCAL2_DX_LOOP_RST_CFG       ),
.RXCKCAL2_D_LOOP_RST_CFG       (RXCKCAL2_D_LOOP_RST_CFG        ),
.RXCKCAL2_S_LOOP_RST_CFG       (RXCKCAL2_S_LOOP_RST_CFG        ),
.RXCKCAL2_X_LOOP_RST_CFG       (RXCKCAL2_X_LOOP_RST_CFG        ),
.RXDFELPMRESET_TIME            (RXDFELPMRESET_TIME             ),
.RXDFELPM_KL_CFG0              (RXDFELPM_KL_CFG0               ),
.RXDFELPM_KL_CFG1              (RXDFELPM_KL_CFG1               ),
.RXDFELPM_KL_CFG2              (RXDFELPM_KL_CFG2               ),
.RXDFE_CFG0                    (RXDFE_CFG0                     ),
.RXDFE_CFG1                    (RXDFE_CFG1                     ),
.RXDFE_GC_CFG0                 (RXDFE_GC_CFG0                  ),
.RXDFE_GC_CFG1                 (RXDFE_GC_CFG1                  ),
.RXDFE_GC_CFG2                 (RXDFE_GC_CFG2                  ),
.RXDFE_H2_CFG0                 (RXDFE_H2_CFG0                  ),
.RXDFE_H2_CFG1                 (RXDFE_H2_CFG1                  ),
.RXDFE_H3_CFG0                 (RXDFE_H3_CFG0                  ),
.RXDFE_H3_CFG1                 (RXDFE_H3_CFG1                  ),
.RXDFE_H4_CFG0                 (RXDFE_H4_CFG0                  ),
.RXDFE_H4_CFG1                 (RXDFE_H4_CFG1                  ),
.RXDFE_H5_CFG0                 (RXDFE_H5_CFG0                  ),
.RXDFE_H5_CFG1                 (RXDFE_H5_CFG1                  ),
.RXDFE_H6_CFG0                 (RXDFE_H6_CFG0                  ),
.RXDFE_H6_CFG1                 (RXDFE_H6_CFG1                  ),
.RXDFE_H7_CFG0                 (RXDFE_H7_CFG0                  ),
.RXDFE_H7_CFG1                 (RXDFE_H7_CFG1                  ),
.RXDFE_H8_CFG0                 (RXDFE_H8_CFG0                  ),
.RXDFE_H8_CFG1                 (RXDFE_H8_CFG1                  ),
.RXDFE_H9_CFG0                 (RXDFE_H9_CFG0                  ),
.RXDFE_H9_CFG1                 (RXDFE_H9_CFG1                  ),
.RXDFE_HA_CFG0                 (RXDFE_HA_CFG0                  ),
.RXDFE_HA_CFG1                 (RXDFE_HA_CFG1                  ),
.RXDFE_HB_CFG0                 (RXDFE_HB_CFG0                  ),
.RXDFE_HB_CFG1                 (RXDFE_HB_CFG1                  ),
.RXDFE_HC_CFG0                 (RXDFE_HC_CFG0                  ),
.RXDFE_HC_CFG1                 (RXDFE_HC_CFG1                  ),
.RXDFE_HD_CFG0                 (RXDFE_HD_CFG0                  ),
.RXDFE_HD_CFG1                 (RXDFE_HD_CFG1                  ),
.RXDFE_HE_CFG0                 (RXDFE_HE_CFG0                  ),
.RXDFE_HE_CFG1                 (RXDFE_HE_CFG1                  ),
.RXDFE_HF_CFG0                 (RXDFE_HF_CFG0                  ),
.RXDFE_HF_CFG1                 (RXDFE_HF_CFG1                  ),
.RXDFE_KH_CFG0                 (RXDFE_KH_CFG0                  ),
.RXDFE_KH_CFG1                 (RXDFE_KH_CFG1                  ),
.RXDFE_KH_CFG2                 (RXDFE_KH_CFG2                  ),
.RXDFE_KH_CFG3                 (RXDFE_KH_CFG3                  ),
.RXDFE_OS_CFG0                 (RXDFE_OS_CFG0                  ),
.RXDFE_OS_CFG1                 (RXDFE_OS_CFG1                  ),
.RXDFE_UT_CFG0                 (RXDFE_UT_CFG0                  ),
.RXDFE_UT_CFG1                 (RXDFE_UT_CFG1                  ),
.RXDFE_UT_CFG2                 (RXDFE_UT_CFG2                  ),
.RXDFE_VP_CFG0                 (RXDFE_VP_CFG0                  ),
.RXDFE_VP_CFG1                 (RXDFE_VP_CFG1                  ),
.RXDLY_CFG                     (RXDLY_CFG                      ),
.RXDLY_LCFG                    (RXDLY_LCFG                     ),
.RXDLY_RAW_CFG                 (RXDLY_RAW_CFG                  ),
.RXDLY_RAW_LCFG                (RXDLY_RAW_LCFG                 ),
.RXELECIDLE_CFG                (RXELECIDLE_CFG                 ),
.RXGBOX_FIFO_INIT_RD_ADDR      (RXGBOX_FIFO_INIT_RD_ADDR       ),
.RXGEARBOX_EN                  (RXGEARBOX_EN                   ),
.RXISCANRESET_TIME             (RXISCANRESET_TIME              ),
.RXLPM_CFG                     (RXLPM_CFG                      ),
.RXLPM_GC_CFG                  (RXLPM_GC_CFG                   ),
.RXLPM_KH_CFG0                 (RXLPM_KH_CFG0                  ),
.RXLPM_KH_CFG1                 (RXLPM_KH_CFG1                  ),
.RXLPM_OS_CFG0                 (RXLPM_OS_CFG0                  ),
.RXLPM_OS_CFG1                 (RXLPM_OS_CFG1                  ),
.RXOSCALRESET_TIME             (RXOSCALRESET_TIME              ),
.RXOUT_DIV                     (RXOUT_DIV                      ),
.RXPCSRESET_TIME               (RXPCSRESET_TIME                ),
.RXPHBEACON_CFG                (RXPHBEACON_CFG                 ),
.RXPHBEACON_RAW_CFG            (RXPHBEACON_RAW_CFG             ),
.RXPHDLY_CFG                   (RXPHDLY_CFG                    ),
.RXPHSAMP_CFG                  (RXPHSAMP_CFG                   ),
.RXPHSAMP_RAW_CFG              (RXPHSAMP_RAW_CFG               ),
.RXPHSLIP_CFG                  (RXPHSLIP_CFG                   ),
.RXPHSLIP_RAW_CFG              (RXPHSLIP_RAW_CFG               ),
.RXPH_MONITOR_SEL              (RXPH_MONITOR_SEL               ),
.RXPI_CFG0                     (RXPI_CFG0                      ),
.RXPI_CFG1                     (RXPI_CFG1                      ),
.RXPMACLK_SEL                  (RXPMACLK_SEL                   ),
.RXPMARESET_TIME               (RXPMARESET_TIME                ),
.RXPRBS_ERR_LOOPBACK           (RXPRBS_ERR_LOOPBACK            ),
.RXPRBS_LINKACQ_CNT            (RXPRBS_LINKACQ_CNT             ),
.RXREFCLKDIV2_SEL              (RXREFCLKDIV2_SEL               ),
.RXSLIDE_AUTO_WAIT             (RXSLIDE_AUTO_WAIT              ),
.RXSLIDE_MODE                  (RXSLIDE_MODE                   ),
.RXSYNC_MULTILANE              (RXSYNC_MULTILANE               ),
.RXSYNC_OVRD                   (RXSYNC_OVRD                    ),
.RXSYNC_SKIP_DA                (RXSYNC_SKIP_DA                 ),
.RX_AFE_CM_EN                  (RX_AFE_CM_EN                   ),
.RX_BIAS_CFG0                  (RX_BIAS_CFG0                   ),
.RX_CAPFF_SARC_ENB             (RX_CAPFF_SARC_ENB              ),
.RX_CLK25_DIV                  (RX_CLK25_DIV                   ),
.RX_CLKMUX_EN                  (RX_CLKMUX_EN                   ),
.RX_CLK_SLIP_OVRD              (RX_CLK_SLIP_OVRD               ),
.RX_CM_BUF_CFG                 (RX_CM_BUF_CFG                  ),
.RX_CM_BUF_PD                  (RX_CM_BUF_PD                   ),
.RX_CM_SEL                     (RX_CM_SEL                      ),
.RX_CM_TRIM                    (RX_CM_TRIM                     ),
.RX_CTLE_PWR_SAVING            (RX_CTLE_PWR_SAVING             ),
.RX_CTLE_RES_CTRL              (RX_CTLE_RES_CTRL               ),
.RX_DATA_WIDTH                 (RX_DATA_WIDTH                  ),
.RX_DDI_SEL                    (RX_DDI_SEL                     ),
.RX_DEGEN_CTRL                 (RX_DEGEN_CTRL                  ),
.RX_DFELPM_CFG0                (RX_DFELPM_CFG0                 ),
.RX_DFELPM_CFG1                (RX_DFELPM_CFG1                 ),
.RX_DFELPM_KLKH_AGC_STUP_EN    (RX_DFELPM_KLKH_AGC_STUP_EN     ),
.RX_DFE_AGC_CFG1               (RX_DFE_AGC_CFG1                ),
.RX_DFE_KL_LPM_KH_CFG0         (RX_DFE_KL_LPM_KH_CFG0          ),
.RX_DFE_KL_LPM_KH_CFG1         (RX_DFE_KL_LPM_KH_CFG1          ),
.RX_DFE_KL_LPM_KL_CFG0         (RX_DFE_KL_LPM_KL_CFG0          ),
.RX_DFE_KL_LPM_KL_CFG1         (RX_DFE_KL_LPM_KL_CFG1          ),
.RX_DFE_LPM_HOLD_DURING_EIDLE  (RX_DFE_LPM_HOLD_DURING_EIDLE   ),
.RX_DISPERR_SEQ_MATCH          (RX_DISPERR_SEQ_MATCH           ),
.RX_DIVRESET_TIME              (RX_DIVRESET_TIME               ),
.RX_EN_CTLE_RCAL_B             (RX_EN_CTLE_RCAL_B              ),
.RX_EN_SUM_RCAL_B              (RX_EN_SUM_RCAL_B               ),
.RX_EYESCAN_VS_CODE            (RX_EYESCAN_VS_CODE             ),
.RX_EYESCAN_VS_NEG_DIR         (RX_EYESCAN_VS_NEG_DIR          ),
.RX_EYESCAN_VS_RANGE           (RX_EYESCAN_VS_RANGE            ),
.RX_EYESCAN_VS_UT_SIGN         (RX_EYESCAN_VS_UT_SIGN          ),
.RX_I2V_FILTER_EN              (RX_I2V_FILTER_EN               ),
.RX_INT_DATAWIDTH              (RX_INT_DATAWIDTH               ),
.RX_PMA_POWER_SAVE             (RX_PMA_POWER_SAVE              ),
.RX_PMA_RSV0                   (RX_PMA_RSV0                    ),
.RX_PROGDIV_CFG                (RX_PROGDIV_CFG                 ),
.RX_PROGDIV_RATE               (RX_PROGDIV_RATE                ),
.RX_RESLOAD_CTRL               (RX_RESLOAD_CTRL                ),
.RX_RESLOAD_OVRD               (RX_RESLOAD_OVRD                ),
.RX_SAMPLE_PERIOD              (RX_SAMPLE_PERIOD               ),
.RX_SIG_VALID_DLY              (RX_SIG_VALID_DLY               ),
.RX_SUM_DEGEN_AVTT_OVERITE     (RX_SUM_DEGEN_AVTT_OVERITE      ),
.RX_SUM_DFETAPREP_EN           (RX_SUM_DFETAPREP_EN            ),
.RX_SUM_IREF_TUNE              (RX_SUM_IREF_TUNE               ),
.RX_SUM_PWR_SAVING             (RX_SUM_PWR_SAVING              ),
.RX_SUM_RES_CTRL               (RX_SUM_RES_CTRL                ),
.RX_SUM_VCMTUNE                (RX_SUM_VCMTUNE                 ),
.RX_SUM_VCM_BIAS_TUNE_EN       (RX_SUM_VCM_BIAS_TUNE_EN        ),
.RX_SUM_VCM_OVWR               (RX_SUM_VCM_OVWR                ),
.RX_SUM_VREF_TUNE              (RX_SUM_VREF_TUNE               ),
.RX_TUNE_AFE_OS                (RX_TUNE_AFE_OS                 ),
.RX_VREG_CTRL                  (RX_VREG_CTRL                   ),
.RX_VREG_PDB                   (RX_VREG_PDB                    ),
.RX_WIDEMODE_CDR               (RX_WIDEMODE_CDR                ),
.RX_WIDEMODE_CDR_GEN3          (RX_WIDEMODE_CDR_GEN3           ),
.RX_WIDEMODE_CDR_GEN4          (RX_WIDEMODE_CDR_GEN4           ),
.RX_XCLK_SEL                   (RX_XCLK_SEL                    ),
.RX_XMODE_SEL                  (RX_XMODE_SEL                   ),
.SAMPLE_CLK_PHASE              (SAMPLE_CLK_PHASE               ),
.SATA_CPLL_CFG                 (SATA_CPLL_CFG                  ),
.SIM_MODE                      (SIM_MODE                       ),
.SIM_RESET_SPEEDUP             (SIM_RESET_SPEEDUP              ),
.SIM_TX_EIDLE_DRIVE_LEVEL      (SIM_TX_EIDLE_DRIVE_LEVEL       ),
.SRSTMODE                      (SRSTMODE                       ),
.TAPDLY_SET_TX                 (TAPDLY_SET_TX                  ),
.TCO_NEW_CFG0                  (TCO_NEW_CFG0                   ),
.TCO_NEW_CFG1                  (TCO_NEW_CFG1                   ),
.TCO_NEW_CFG2                  (TCO_NEW_CFG2                   ),
.TCO_NEW_CFG3                  (TCO_NEW_CFG3                   ),
.TCO_RSVD1                     (TCO_RSVD1                      ),
.TCO_RSVD2                     (TCO_RSVD2                      ),
.TERM_RCAL_CFG                 (TERM_RCAL_CFG                  ),
.TERM_RCAL_OVRD                (TERM_RCAL_OVRD                 ),
.TRANS_TIME_RATE               (TRANS_TIME_RATE                ),
.TST_RSV0                      (TST_RSV0                       ),
.TST_RSV1                      (TST_RSV1                       ),
.TXBUF_EN                      (TXBUF_EN                       ),
.TXDLY_CFG                     (TXDLY_CFG                      ),
.TXDLY_LCFG                    (TXDLY_LCFG                     ),
.TXDRV_FREQBAND                (TXDRV_FREQBAND                 ),
.TXFE_CFG0                     (TXFE_CFG0                      ),
.TXFE_CFG1                     (TXFE_CFG1                      ),
.TXFE_CFG2                     (TXFE_CFG2                      ),
.TXFE_CFG3                     (TXFE_CFG3                      ),
.TXFIFO_ADDR_CFG               (TXFIFO_ADDR_CFG                ),
.TXGBOX_FIFO_INIT_RD_ADDR      (TXGBOX_FIFO_INIT_RD_ADDR       ),
.TXOUT_DIV                     (TXOUT_DIV                      ),
.TXPCSRESET_TIME               (TXPCSRESET_TIME                ),
.TXPHDLY_CFG0                  (TXPHDLY_CFG0                   ),
.TXPHDLY_CFG1                  (TXPHDLY_CFG1                   ),
.TXPH_CFG                      (TXPH_CFG                       ),
.TXPH_CFG2                     (TXPH_CFG2                      ),
.TXPH_MONITOR_SEL              (TXPH_MONITOR_SEL               ),
.TXPI_CFG0                     (TXPI_CFG0                      ),
.TXPI_CFG1                     (TXPI_CFG1                      ),
.TXPI_GRAY_SEL                 (TXPI_GRAY_SEL                  ),
.TXPI_INVSTROBE_SEL            (TXPI_INVSTROBE_SEL             ),
.TXPI_PPM                      (TXPI_PPM                       ),
.TXPI_PPM_CFG                  (TXPI_PPM_CFG                   ),
.TXPI_SYNFREQ_PPM              (TXPI_SYNFREQ_PPM               ),
.TXPMARESET_TIME               (TXPMARESET_TIME                ),
.TXREFCLKDIV2_SEL              (TXREFCLKDIV2_SEL               ),
.TXSWBST_BST                   (TXSWBST_BST                    ),
.TXSWBST_EN                    (TXSWBST_EN                     ),
.TXSWBST_MAG                   (TXSWBST_MAG                    ),
.TXSYNC_MULTILANE              (TXSYNC_MULTILANE               ),
.TXSYNC_OVRD                   (TXSYNC_OVRD                    ),
.TXSYNC_SKIP_DA                (TXSYNC_SKIP_DA                 ),
.TX_CLK25_DIV                  (TX_CLK25_DIV                   ),
.TX_CLKMUX_EN                  (TX_CLKMUX_EN                   ),
.TX_DATA_WIDTH                 (TX_DATA_WIDTH                  ),
.TX_DCC_LOOP_RST_CFG           (TX_DCC_LOOP_RST_CFG            ),
.TX_DIVRESET_TIME              (TX_DIVRESET_TIME               ),
.TX_EIDLE_ASSERT_DELAY         (TX_EIDLE_ASSERT_DELAY          ),
.TX_EIDLE_DEASSERT_DELAY       (TX_EIDLE_DEASSERT_DELAY        ),
.TX_FABINT_USRCLK_FLOP         (TX_FABINT_USRCLK_FLOP          ),
.TX_FIFO_BYP_EN                (TX_FIFO_BYP_EN                 ),
.TX_IDLE_DATA_ZERO             (TX_IDLE_DATA_ZERO              ),
.TX_INT_DATAWIDTH              (TX_INT_DATAWIDTH               ),
.TX_LOOPBACK_DRIVE_HIZ         (TX_LOOPBACK_DRIVE_HIZ          ),
.TX_MAINCURSOR_SEL             (TX_MAINCURSOR_SEL              ),
.TX_PHICAL_CFG0                (TX_PHICAL_CFG0                 ),
.TX_PHICAL_CFG1                (TX_PHICAL_CFG1                 ),
.TX_PI_BIASSET                 (TX_PI_BIASSET                  ),
.TX_PMADATA_OPT                (TX_PMADATA_OPT                 ),
.TX_PMA_POWER_SAVE             (TX_PMA_POWER_SAVE              ),
.TX_PMA_RSV0                   (TX_PMA_RSV0                    ),
.TX_PMA_RSV1                   (TX_PMA_RSV1                    ),
.TX_PROGCLK_SEL                (TX_PROGCLK_SEL                 ),
.TX_PROGDIV_CFG                (TX_PROGDIV_CFG                 ),
.TX_PROGDIV_RATE               (TX_PROGDIV_RATE                ),
.TX_SAMPLE_PERIOD              (TX_SAMPLE_PERIOD               ),
.TX_SW_MEAS                    (TX_SW_MEAS                     ),
.TX_VREG_CTRL                  (TX_VREG_CTRL                   ),
.TX_VREG_PDB                   (TX_VREG_PDB                    ),
.TX_VREG_VREFSEL               (TX_VREG_VREFSEL                ),
.TX_XCLK_SEL                   (TX_XCLK_SEL                    ),
.USE_PCS_CLK_PHASE_SEL         (USE_PCS_CLK_PHASE_SEL          ),
.USE_RAW_ELEC                  (USE_RAW_ELEC                   ),
.Y_ALL_MODE                    (Y_ALL_MODE                     )
) gtf_channel_inst (
 .CDRSTEPDIR                (gtf_ch_cdrstepdir                ),
 .CDRSTEPSQ                 (gtf_ch_cdrstepsq                 ),
 .CDRSTEPSX                 (gtf_ch_cdrstepsx                 ),
 .CFGRESET                  (gtf_ch_cfgreset                  ),
 .CLKRSVD0                  (gtf_ch_clkrsvd0                  ),
 .CLKRSVD1                  (gtf_ch_clkrsvd1                  ),
 .CPLLFREQLOCK              (gtf_ch_cpllfreqlock              ),
 .CPLLLOCKDETCLK            (gtf_ch_cplllockdetclk            ),
 .CPLLLOCKEN                (gtf_ch_cplllocken                ),
 .CPLLPD                    (gtf_ch_cpllpd                    ),
 .CPLLRESET                 (gtf_ch_cpllreset                 ),
 .CTLTXRESENDPAUSE          (gtf_ch_ctltxresendpause          ),
 .CTLTXSENDIDLE             (gtf_ch_ctltxsendidle             ),
 .CTLTXSENDLFI              (gtf_ch_ctltxsendlfi              ),
 .CTLTXSENDRFI              (gtf_ch_ctltxsendrfi              ),
 .DMONFIFORESET             (gtf_ch_dmonfiforeset             ),
 .DMONITORCLK               (gtf_ch_dmonitorclk               ),
 .DRPCLK                    (gtf_ch_drpclk                    ),
 .DRPEN                     (gtf_ch_drpen                     ),
 .DRPRST                    (gtf_ch_drprst                    ),
 .DRPWE                     (gtf_ch_drpwe                     ),
 .EYESCANRESET              (gtf_ch_eyescanreset              ),
 .EYESCANTRIGGER            (gtf_ch_eyescantrigger            ),
 .FREQOS                    (gtf_ch_freqos                    ),
 .GTFRXN                    (gtf_ch_gtfrxn                    ),
 .GTFRXP                    (gtf_ch_gtfrxp                    ),
 .GTGREFCLK                 (gtf_ch_gtgrefclk                 ),
 .GTNORTHREFCLK0            (gtf_ch_gtnorthrefclk0            ),
 .GTNORTHREFCLK1            (gtf_ch_gtnorthrefclk1            ),
 .GTREFCLK0                 (gtf_ch_gtrefclk0                 ),
 .GTREFCLK1                 (gtf_ch_gtrefclk1                 ),
 .GTRXRESET                 (gtf_ch_gtrxreset                 ),
 .GTRXRESETSEL              (gtf_ch_gtrxresetsel              ),
 .GTSOUTHREFCLK0            (gtf_ch_gtsouthrefclk0            ),
 .GTSOUTHREFCLK1            (gtf_ch_gtsouthrefclk1            ),
 .GTTXRESET                 (gtf_ch_gttxreset                 ),
 .GTTXRESETSEL              (gtf_ch_gttxresetsel              ),
 .INCPCTRL                  (gtf_ch_incpctrl                  ),
 .QPLL0CLK                  (gtf_ch_qpll0clk                  ),
 .QPLL0FREQLOCK             (gtf_ch_qpll0freqlock             ),
 .QPLL0REFCLK               (gtf_ch_qpll0refclk               ),
 .QPLL1CLK                  (gtf_ch_qpll1clk                  ),
 .QPLL1FREQLOCK             (gtf_ch_qpll1freqlock             ),
 .QPLL1REFCLK               (gtf_ch_qpll1refclk               ),
 .RESETOVRD                 (gtf_ch_resetovrd                 ),
 .RXAFECFOKEN               (gtf_ch_rxafecfoken               ),
 .RXCDRFREQRESET            (gtf_ch_rxcdrfreqreset            ),
 .RXCDRHOLD                 (gtf_ch_rxcdrhold                 ),
 .RXCDROVRDEN               (gtf_ch_rxcdrovrden               ),
 .RXCDRRESET                (gtf_ch_rxcdrreset                ),
 .RXCKCALRESET              (gtf_ch_rxckcalreset              ),
 .RXDFEAGCHOLD              (gtf_ch_rxdfeagchold              ),
 .RXDFEAGCOVRDEN            (gtf_ch_rxdfeagcovrden            ),
 .RXDFECFOKFEN              (gtf_ch_rxdfecfokfen              ),
 .RXDFECFOKFPULSE           (gtf_ch_rxdfecfokfpulse           ),
 .RXDFECFOKHOLD             (gtf_ch_rxdfecfokhold             ),
 .RXDFECFOKOVREN            (gtf_ch_rxdfecfokovren            ),
 .RXDFEKHHOLD               (gtf_ch_rxdfekhhold               ),
 .RXDFEKHOVRDEN             (gtf_ch_rxdfekhovrden             ),
 .RXDFELFHOLD               (gtf_ch_rxdfelfhold               ),
 .RXDFELFOVRDEN             (gtf_ch_rxdfelfovrden             ),
 .RXDFELPMRESET             (gtf_ch_rxdfelpmreset             ),
 .RXDFETAP10HOLD            (gtf_ch_rxdfetap10hold            ),
 .RXDFETAP10OVRDEN          (gtf_ch_rxdfetap10ovrden          ),
 .RXDFETAP11HOLD            (gtf_ch_rxdfetap11hold            ),
 .RXDFETAP11OVRDEN          (gtf_ch_rxdfetap11ovrden          ),
 .RXDFETAP12HOLD            (gtf_ch_rxdfetap12hold            ),
 .RXDFETAP12OVRDEN          (gtf_ch_rxdfetap12ovrden          ),
 .RXDFETAP13HOLD            (gtf_ch_rxdfetap13hold            ),
 .RXDFETAP13OVRDEN          (gtf_ch_rxdfetap13ovrden          ),
 .RXDFETAP14HOLD            (gtf_ch_rxdfetap14hold            ),
 .RXDFETAP14OVRDEN          (gtf_ch_rxdfetap14ovrden          ),
 .RXDFETAP15HOLD            (gtf_ch_rxdfetap15hold            ),
 .RXDFETAP15OVRDEN          (gtf_ch_rxdfetap15ovrden          ),
 .RXDFETAP2HOLD             (gtf_ch_rxdfetap2hold             ),
 .RXDFETAP2OVRDEN           (gtf_ch_rxdfetap2ovrden           ),
 .RXDFETAP3HOLD             (gtf_ch_rxdfetap3hold             ),
 .RXDFETAP3OVRDEN           (gtf_ch_rxdfetap3ovrden           ),
 .RXDFETAP4HOLD             (gtf_ch_rxdfetap4hold             ),
 .RXDFETAP4OVRDEN           (gtf_ch_rxdfetap4ovrden           ),
 .RXDFETAP5HOLD             (gtf_ch_rxdfetap5hold             ),
 .RXDFETAP5OVRDEN           (gtf_ch_rxdfetap5ovrden           ),
 .RXDFETAP6HOLD             (gtf_ch_rxdfetap6hold             ),
 .RXDFETAP6OVRDEN           (gtf_ch_rxdfetap6ovrden           ),
 .RXDFETAP7HOLD             (gtf_ch_rxdfetap7hold             ),
 .RXDFETAP7OVRDEN           (gtf_ch_rxdfetap7ovrden           ),
 .RXDFETAP8HOLD             (gtf_ch_rxdfetap8hold             ),
 .RXDFETAP8OVRDEN           (gtf_ch_rxdfetap8ovrden           ),
 .RXDFETAP9HOLD             (gtf_ch_rxdfetap9hold             ),
 .RXDFETAP9OVRDEN           (gtf_ch_rxdfetap9ovrden           ),
 .RXDFEUTHOLD               (gtf_ch_rxdfeuthold               ),
 .RXDFEUTOVRDEN             (gtf_ch_rxdfeutovrden             ),
 .RXDFEVPHOLD               (gtf_ch_rxdfevphold               ),
 .RXDFEVPOVRDEN             (gtf_ch_rxdfevpovrden             ),
 .RXDFEXYDEN                (gtf_ch_rxdfexyden                ),
 .RXDLYBYPASS               (gtf_ch_rxdlybypass               ),
 .RXDLYEN                   (gtf_ch_rxdlyen                   ),
 .RXDLYOVRDEN               (gtf_ch_rxdlyovrden               ),
 .RXDLYSRESET               (gtf_ch_rxdlysreset               ),
 .RXLPMEN                   (gtf_ch_rxlpmen                   ),
 .RXLPMGCHOLD               (gtf_ch_rxlpmgchold               ),
 .RXLPMGCOVRDEN             (gtf_ch_rxlpmgcovrden             ),
 .RXLPMHFHOLD               (gtf_ch_rxlpmhfhold               ),
 .RXLPMHFOVRDEN             (gtf_ch_rxlpmhfovrden             ),
 .RXLPMLFHOLD               (gtf_ch_rxlpmlfhold               ),
 .RXLPMLFKLOVRDEN           (gtf_ch_rxlpmlfklovrden           ),
 .RXLPMOSHOLD               (gtf_ch_rxlpmoshold               ),
 .RXLPMOSOVRDEN             (gtf_ch_rxlpmosovrden             ),
 .RXOSCALRESET              (gtf_ch_rxoscalreset              ),
 .RXOSHOLD                  (gtf_ch_rxoshold                  ),
 .RXOSOVRDEN                (gtf_ch_rxosovrden                ),
 .RXPCSRESET                (gtf_ch_rxpcsreset                ),
 .RXPHALIGN                 (gtf_ch_rxphalign                 ),
 .RXPHALIGNEN               (gtf_ch_rxphalignen               ),
 .RXPHDLYPD                 (gtf_ch_rxphdlypd                 ),
 .RXPHDLYRESET              (gtf_ch_rxphdlyreset              ),
 .RXPMARESET                (gtf_ch_rxpmareset                ),
 .RXPOLARITY                (gtf_ch_rxpolarity                ),
 .RXPRBSCNTRESET            (gtf_ch_rxprbscntreset            ),
 .RXPROGDIVRESET            (gtf_ch_rxprogdivreset            ),
 .RXSLIPOUTCLK              (gtf_ch_rxslipoutclk              ),
 .RXSLIPPMA                 (gtf_ch_rxslippma                 ),
 .RXSYNCALLIN               (gtf_ch_rxsyncallin               ),
 .RXSYNCIN                  (gtf_ch_rxsyncin                  ),
 .RXSYNCMODE                (gtf_ch_rxsyncmode                ),
 .RXTERMINATION             (gtf_ch_rxtermination             ),
 .RXUSERRDY                 (gtf_ch_rxuserrdy                 ),
 .RXUSRCLK                  (gtf_ch_rxusrclk                  ),
 .RXUSRCLK2                 (gtf_ch_rxusrclk2                 ),
 .TXAXISTERR                (gtf_ch_txaxisterr                ),
 .TXAXISTPOISON             (gtf_ch_txaxistpoison             ),
 .TXAXISTVALID              (gtf_ch_txaxistvalid              ),
 .TXDCCFORCESTART           (gtf_ch_txdccforcestart           ),
 .TXDCCRESET                (gtf_ch_txdccreset                ),
 .TXDLYBYPASS               (gtf_ch_txdlybypass               ),
 .TXDLYEN                   (gtf_ch_txdlyen                   ),
 .TXDLYHOLD                 (gtf_ch_txdlyhold                 ),
 .TXDLYOVRDEN               (gtf_ch_txdlyovrden               ),
 .TXDLYSRESET               (gtf_ch_txdlysreset               ),
 .TXDLYUPDOWN               (gtf_ch_txdlyupdown               ),
 .TXELECIDLE                (gtf_ch_txelecidle                ),
 .TXGBSEQSYNC               (gtf_ch_txgbseqsync               ),
 .TXMUXDCDEXHOLD            (gtf_ch_txmuxdcdexhold            ),
 .TXMUXDCDORWREN            (gtf_ch_txmuxdcdorwren            ),
 .TXPCSRESET                (gtf_ch_txpcsreset                ),
 .TXPHALIGN                 (gtf_ch_txphalign                 ),
 .TXPHALIGNEN               (gtf_ch_txphalignen               ),
 .TXPHDLYPD                 (gtf_ch_txphdlypd                 ),
 .TXPHDLYRESET              (gtf_ch_txphdlyreset              ),
 .TXPHDLYTSTCLK             (gtf_ch_txphdlytstclk             ),
 .TXPHINIT                  (gtf_ch_txphinit                  ),
 .TXPHOVRDEN                (gtf_ch_txphovrden                ),
 .TXPIPPMEN                 (gtf_ch_txpippmen                 ),
 .TXPIPPMOVRDEN             (gtf_ch_txpippmovrden             ),
 .TXPIPPMPD                 (gtf_ch_txpippmpd                 ),
 .TXPIPPMSEL                (gtf_ch_txpippmsel                ),
 .TXPISOPD                  (gtf_ch_txpisopd                  ),
 .TXPMARESET                (gtf_ch_txpmareset                ),
 .TXPOLARITY                (gtf_ch_txpolarity                ),
 .TXPRBSFORCEERR            (gtf_ch_txprbsforceerr            ),
 .TXPROGDIVRESET            (gtf_ch_txprogdivreset            ),
 .TXSYNCALLIN               (gtf_ch_txsyncallin               ),
 .TXSYNCIN                  (gtf_ch_txsyncin                  ),
 .TXSYNCMODE                (gtf_ch_txsyncmode                ),
 .TXUSERRDY                 (gtf_ch_txuserrdy                 ),
 .TXUSRCLK                  (gtf_ch_txusrclk                  ),
 .TXUSRCLK2                 (gtf_ch_txusrclk2                 ),
 .DRPDI                     (gtf_ch_drpdi                     ),
 .GTRSVD                    (gtf_ch_gtrsvd                    ),
 .PCSRSVDIN                 (gtf_ch_pcsrsvdin                 ),
 .TSTIN                     (gtf_ch_tstin                     ),
 .RXELECIDLEMODE            (gtf_ch_rxelecidlemode            ),
 .RXMONITORSEL              (gtf_ch_rxmonitorsel              ),
 .RXPD                      (gtf_ch_rxpd                      ),
 .RXPLLCLKSEL               (gtf_ch_rxpllclksel               ),
 .RXSYSCLKSEL               (gtf_ch_rxsysclksel               ),
 .TXAXISTSOF                (gtf_ch_txaxistsof                ),
 .TXPD                      (gtf_ch_txpd                      ),
 .TXPLLCLKSEL               (gtf_ch_txpllclksel               ),
 .TXSYSCLKSEL               (gtf_ch_txsysclksel               ),
 .CPLLREFCLKSEL             (gtf_ch_cpllrefclksel             ),
 .LOOPBACK                  (gtf_ch_loopback                  ),
 .RXOUTCLKSEL               (gtf_ch_rxoutclksel               ),
 .TXOUTCLKSEL               (gtf_ch_txoutclksel               ),
 .TXRAWDATA                 (gtf_ch_txrawdata                 ),
 .RXDFECFOKFCNUM            (gtf_ch_rxdfecfokfcnum            ),
 .RXPRBSSEL                 (gtf_ch_rxprbssel                 ),
 .TXPRBSSEL                 (gtf_ch_txprbssel                 ),
 .TXAXISTTERM               (gtf_ch_txaxistterm               ),
 .TXDIFFCTRL                (gtf_ch_txdiffctrl                ),
 .TXPIPPMSTEPSIZE           (gtf_ch_txpippmstepsize           ),
 .TXPOSTCURSOR              (gtf_ch_txpostcursor              ),
 .TXPRECURSOR               (gtf_ch_txprecursor               ),
 .TXAXISTDATA               (gtf_ch_txaxistdata               ),
 .RXCKCALSTART              (gtf_ch_rxckcalstart              ),
 .TXMAINCURSOR              (gtf_ch_txmaincursor              ),
 .TXAXISTLAST               (gtf_ch_txaxistlast               ),
 .TXAXISTPRE                (gtf_ch_txaxistpre                ),
 .CTLRXPAUSEACK             (gtf_ch_ctlrxpauseack             ),
 .CTLTXPAUSEREQ             (gtf_ch_ctltxpausereq             ),
 .DRPADDR                   (gtf_ch_drpaddr                   ),
 .CPLLFBCLKLOST             (gtf_ch_cpllfbclklost             ),
 .CPLLLOCK                  (gtf_ch_cplllock                  ),
 .CPLLREFCLKLOST            (gtf_ch_cpllrefclklost            ),
 .DMONITOROUTCLK            (gtf_ch_dmonitoroutclk            ),
 .DRPRDY                    (gtf_ch_drprdy                    ),
 .EYESCANDATAERROR          (gtf_ch_eyescandataerror          ),
 .GTFTXN                    (gtf_ch_gtftxn                    ),
 .GTFTXP                    (gtf_ch_gtftxp                    ),
 .GTPOWERGOOD               (gtf_ch_gtpowergood               ),
 .GTREFCLKMONITOR           (gtf_ch_gtrefclkmonitor           ),
 .RESETEXCEPTION            (gtf_ch_resetexception            ),
 .RXAXISTERR                (gtf_ch_rxaxisterr                ),
 .RXAXISTVALID              (gtf_ch_rxaxistvalid              ),
 .RXBITSLIP                 (gtf_ch_rxbitslip                 ),
 .RXCDRLOCK                 (gtf_ch_rxcdrlock                 ),
 .RXCDRPHDONE               (gtf_ch_rxcdrphdone               ),
 .RXCKCALDONE               (gtf_ch_rxckcaldone               ),
 .RXDLYSRESETDONE           (gtf_ch_rxdlysresetdone           ),
 .RXELECIDLE                (gtf_ch_rxelecidle                ),
 .RXGBSEQSTART              (gtf_ch_rxgbseqstart              ),
 .RXOSINTDONE               (gtf_ch_rxosintdone               ),
 .RXOSINTSTARTED            (gtf_ch_rxosintstarted            ),
 .RXOSINTSTROBEDONE         (gtf_ch_rxosintstrobedone         ),
 .RXOSINTSTROBESTARTED      (gtf_ch_rxosintstrobestarted      ),
 .RXOUTCLK                  (gtf_ch_rxoutclk                  ),
 .RXOUTCLKFABRIC            (gtf_ch_rxoutclkfabric            ),
 .RXOUTCLKPCS               (gtf_ch_rxoutclkpcs               ),
 .RXPHALIGNDONE             (gtf_ch_rxphaligndone             ),
 .RXPHALIGNERR              (gtf_ch_rxphalignerr              ),
 .RXPMARESETDONE            (gtf_ch_rxpmaresetdone            ),
 .RXPRBSERR                 (gtf_ch_rxprbserr                 ),
 .RXPRBSLOCKED              (gtf_ch_rxprbslocked              ),
 .RXPRGDIVRESETDONE         (gtf_ch_rxprgdivresetdone         ),
 .RXPTPSOP                  (gtf_ch_rxptpsop                  ),
 .RXPTPSOPPOS               (gtf_ch_rxptpsoppos               ),
 .RXRECCLKOUT               (gtf_ch_rxrecclkout               ),
 .RXRESETDONE               (gtf_ch_rxresetdone               ),
 .RXSLIPDONE                (gtf_ch_rxslipdone                ),
 .RXSLIPOUTCLKRDY           (gtf_ch_rxslipoutclkrdy           ),
 .RXSLIPPMARDY              (gtf_ch_rxslippmardy              ),
 .RXSYNCDONE                (gtf_ch_rxsyncdone                ),
 .RXSYNCOUT                 (gtf_ch_rxsyncout                 ),
 .STATRXBADCODE             (gtf_ch_statrxbadcode             ),
 .STATRXBADFCS              (gtf_ch_statrxbadfcs              ),
 .STATRXBADPREAMBLE         (gtf_ch_statrxbadpreamble         ),
 .STATRXBADSFD              (gtf_ch_statrxbadsfd              ),
 .STATRXBLOCKLOCK           (gtf_ch_statrxblocklock           ),
 .STATRXBROADCAST           (gtf_ch_statrxbroadcast           ),
 .STATRXFCSERR              (gtf_ch_statrxfcserr              ),
 .STATRXFRAMINGERR          (gtf_ch_statrxframingerr          ),
 .STATRXGOTSIGNALOS         (gtf_ch_statrxgotsignalos         ),
 .STATRXHIBER               (gtf_ch_statrxhiber               ),
 .STATRXINRANGEERR          (gtf_ch_statrxinrangeerr          ),
 .STATRXINTERNALLOCALFAULT  (gtf_ch_statrxinternallocalfault  ),
 .STATRXLOCALFAULT          (gtf_ch_statrxlocalfault          ),
 .STATRXMULTICAST           (gtf_ch_statrxmulticast           ),
 .STATRXPKT                 (gtf_ch_statrxpkt                 ),
 .STATRXPKTERR              (gtf_ch_statrxpkterr              ),
 .STATRXRECEIVEDLOCALFAULT  (gtf_ch_statrxreceivedlocalfault  ),
 .STATRXREMOTEFAULT         (gtf_ch_statrxremotefault         ),
 .STATRXSTATUS              (gtf_ch_statrxstatus              ),
 .STATRXSTOMPEDFCS          (gtf_ch_statrxstompedfcs          ),
 .STATRXTESTPATTERNMISMATCH (gtf_ch_statrxtestpatternmismatch ),
 .STATRXTRUNCATED           (gtf_ch_statrxtruncated           ),
 .STATRXUNICAST             (gtf_ch_statrxunicast             ),
 .STATRXVALIDCTRLCODE       (gtf_ch_statrxvalidctrlcode       ),
 .STATRXVLAN                (gtf_ch_statrxvlan                ),
 .STATTXBADFCS              (gtf_ch_stattxbadfcs              ),
 .STATTXBROADCAST           (gtf_ch_stattxbroadcast           ),
 .STATTXFCSERR              (gtf_ch_stattxfcserr              ),
 .STATTXMULTICAST           (gtf_ch_stattxmulticast           ),
 .STATTXPKT                 (gtf_ch_stattxpkt                 ),
 .STATTXPKTERR              (gtf_ch_stattxpkterr              ),
 .STATTXUNICAST             (gtf_ch_stattxunicast             ),
 .STATTXVLAN                (gtf_ch_stattxvlan                ),
 .TXAXISTREADY              (gtf_ch_txaxistready              ),
 .TXDCCDONE                 (gtf_ch_txdccdone                 ),
 .TXDLYSRESETDONE           (gtf_ch_txdlysresetdone           ),
 .TXGBSEQSTART              (gtf_ch_txgbseqstart              ),
 .TXOUTCLK                  (gtf_ch_txoutclk                  ),
 .TXOUTCLKFABRIC            (gtf_ch_txoutclkfabric            ),
 .TXOUTCLKPCS               (gtf_ch_txoutclkpcs               ),
 .TXPHALIGNDONE             (gtf_ch_txphaligndone             ),
 .TXPHINITDONE              (gtf_ch_txphinitdone              ),
 .TXPMARESETDONE            (gtf_ch_txpmaresetdone            ),
 .TXPRGDIVRESETDONE         (gtf_ch_txprgdivresetdone         ),
 .TXPTPSOP                  (gtf_ch_txptpsop                  ),
 .TXPTPSOPPOS               (gtf_ch_txptpsoppos               ),
 .TXRESETDONE               (gtf_ch_txresetdone               ),
 .TXSYNCDONE                (gtf_ch_txsyncdone                ),
 .TXSYNCOUT                 (gtf_ch_txsyncout                 ),
 .TXUNFOUT                  (gtf_ch_txunfout                  ),
 .DMONITOROUT               (gtf_ch_dmonitorout               ),
 .DRPDO                     (gtf_ch_drpdo                     ),
 .PCSRSVDOUT                (gtf_ch_pcsrsvdout                ),
 .PINRSRVDAS                (gtf_ch_pinrsrvdas                ),
 .RXAXISTSOF                (gtf_ch_rxaxistsof                ),
 .RXRAWDATA                 (gtf_ch_rxrawdata                 ),
 .STATRXBYTES               (gtf_ch_statrxbytes               ),
 .STATTXBYTES               (gtf_ch_stattxbytes               ),
 .RXAXISTTERM               (gtf_ch_rxaxistterm               ),
 .RXAXISTDATA               (gtf_ch_rxaxistdata               ),
 .RXAXISTLAST               (gtf_ch_rxaxistlast               ),
 .RXAXISTPRE                (gtf_ch_rxaxistpre                ),
 .RXMONITOROUT              (gtf_ch_rxmonitorout              ),
 .STATRXPAUSEQUANTA         (gtf_ch_statrxpausequanta         ),
 .STATRXPAUSEREQ            (gtf_ch_statrxpausereq            ),
 .STATRXPAUSEVALID          (gtf_ch_statrxpausevalid          ),
 .STATTXPAUSEVALID          (gtf_ch_stattxpausevalid          )
);
//----}


endmodule
`default_nettype wire
//------}
