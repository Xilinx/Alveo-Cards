/*
Copyright (c) 2023, Advanced Micro Devices, Inc. All rights reserved.
SPDX-License-Identifier: MIT
*/

//------------------------------------------------------------------------------


//------{
`timescale 1fs/1fs
`default_nettype none
(* DowngradeIPIdentifiedWarnings="yes" *)
module gtfwizard_mac_example_gtf_common # (
  parameter [0:0] AEN_QPLL0_FBDIV = 1'b1,
  parameter [0:0] AEN_QPLL1_FBDIV = 1'b1,
  parameter [0:0] AEN_SDM0TOGGLE = 1'b0,
  parameter [0:0] AEN_SDM1TOGGLE = 1'b0,
  parameter [0:0] A_SDM0TOGGLE = 1'b0,
  parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000,
  parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000,
  parameter [0:0] A_SDM1TOGGLE = 1'b0,
  parameter [15:0] BIAS_CFG0 = 16'h0000,
  parameter [15:0] BIAS_CFG1 = 16'h0000,
  parameter [15:0] BIAS_CFG2 = 16'h0000,
  parameter [15:0] BIAS_CFG3 = 16'h0000,
  parameter [15:0] BIAS_CFG4 = 16'h0000,
  parameter [15:0] BIAS_CFG_RSVD = 16'h0000,
  parameter [15:0] COMMON_CFG0 = 16'h0000,
  parameter [15:0] COMMON_CFG1 = 16'h0000,
  parameter [15:0] POR_CFG = 16'h0000,
  parameter [15:0] PPF0_CFG = 16'h0F00,
  parameter [15:0] PPF1_CFG = 16'h0F00,
  parameter QPLL0CLKOUT_RATE = "FULL",
  parameter [15:0] QPLL0_CFG0 = 16'h391C,
  parameter [15:0] QPLL0_CFG1 = 16'h0000,
  parameter [15:0] QPLL0_CFG1_G3 = 16'h0020,
  parameter [15:0] QPLL0_CFG2 = 16'h0F80,
  parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80,
  parameter [15:0] QPLL0_CFG3 = 16'h0120,
  parameter [15:0] QPLL0_CFG4 = 16'h0002,
  parameter [9:0] QPLL0_CP = 10'b0000011111,
  parameter [9:0] QPLL0_CP_G3 = 10'b0000011111,
  parameter integer QPLL0_FBDIV = 66,
  parameter integer QPLL0_FBDIV_G3 = 80,
  parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000,
  parameter [7:0] QPLL0_INIT_CFG1 = 8'h00,
  parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8,
  parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8,
  parameter [9:0] QPLL0_LPF = 10'b1011111111,
  parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111,
  parameter [0:0] QPLL0_PCI_EN = 1'b0,
  parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0,
  parameter integer QPLL0_REFCLK_DIV = 1,
  parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040,
  parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000,
  parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000,
  parameter QPLL1CLKOUT_RATE = "FULL",
  parameter [15:0] QPLL1_CFG0 = 16'h691C,
  parameter [15:0] QPLL1_CFG1 = 16'h0020,
  parameter [15:0] QPLL1_CFG1_G3 = 16'h0020,
  parameter [15:0] QPLL1_CFG2 = 16'h0F80,
  parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80,
  parameter [15:0] QPLL1_CFG3 = 16'h0120,
  parameter [15:0] QPLL1_CFG4 = 16'h0002,
  parameter [9:0] QPLL1_CP = 10'b0000011111,
  parameter [9:0] QPLL1_CP_G3 = 10'b0000011111,
  parameter integer QPLL1_FBDIV = 66,
  parameter integer QPLL1_FBDIV_G3 = 80,
  parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000,
  parameter [7:0] QPLL1_INIT_CFG1 = 8'h00,
  parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8,
  parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8,
  parameter [9:0] QPLL1_LPF = 10'b1011111111,
  parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111,
  parameter [0:0] QPLL1_PCI_EN = 1'b0,
  parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0,
  parameter integer QPLL1_REFCLK_DIV = 1,
  parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000,
  parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000,
  parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000,
  parameter [15:0] RSVD_ATTR0 = 16'h0000,
  parameter [15:0] RSVD_ATTR1 = 16'h0000,
  parameter [15:0] RSVD_ATTR2 = 16'h0000,
  parameter [15:0] RSVD_ATTR3 = 16'h0000,
  parameter [1:0] RXRECCLKOUT0_SEL = 2'b00,
  parameter [1:0] RXRECCLKOUT1_SEL = 2'b00,
  parameter [0:0] SARC_ENB = 1'b0,
  parameter [0:0] SARC_SEL = 1'b0,
  parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000,
  parameter [8:0] SDM0INITSEED0_1 = 9'b000000000,
  parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000,
  parameter [8:0] SDM1INITSEED0_1 = 9'b000000000,
  parameter SIM_MODE = "FAST",
  parameter SIM_RESET_SPEEDUP = "TRUE"
)(
  input  wire         gtf_cm_bgbypassb,
  input  wire         gtf_cm_bgmonitorenb,
  input  wire         gtf_cm_bgpdb,
  input  wire         gtf_cm_bgrcalovrdenb,
  input  wire         gtf_cm_drpclk,
  input  wire         gtf_cm_drpen,
  input  wire         gtf_cm_drpwe,
  input  wire         gtf_cm_gtgrefclk0,
  input  wire         gtf_cm_gtgrefclk1,
  input  wire         gtf_cm_gtnorthrefclk00,
  input  wire         gtf_cm_gtnorthrefclk01,
  input  wire         gtf_cm_gtnorthrefclk10,
  input  wire         gtf_cm_gtnorthrefclk11,
  input  wire         gtf_cm_gtrefclk00,
  input  wire         gtf_cm_gtrefclk01,
  input  wire         gtf_cm_gtrefclk10,
  input  wire         gtf_cm_gtrefclk11,
  input  wire         gtf_cm_gtsouthrefclk00,
  input  wire         gtf_cm_gtsouthrefclk01,
  input  wire         gtf_cm_gtsouthrefclk10,
  input  wire         gtf_cm_gtsouthrefclk11,
  input  wire         gtf_cm_qpll0clkrsvd0,
  input  wire         gtf_cm_qpll0clkrsvd1,
  input  wire         gtf_cm_qpll0lockdetclk,
  input  wire         gtf_cm_qpll0locken,
  input  wire         gtf_cm_qpll0pd,
  input  wire         gtf_cm_qpll0reset,
  input  wire         gtf_cm_qpll1clkrsvd0,
  input  wire         gtf_cm_qpll1clkrsvd1,
  input  wire         gtf_cm_qpll1lockdetclk,
  input  wire         gtf_cm_qpll1locken,
  input  wire         gtf_cm_qpll1pd,
  input  wire         gtf_cm_qpll1reset,
  input  wire         gtf_cm_rcalenb,
  input  wire         gtf_cm_sdm0reset,
  input  wire         gtf_cm_sdm0toggle,
  input  wire         gtf_cm_sdm1reset,
  input  wire         gtf_cm_sdm1toggle,
  input  wire  [15:0] gtf_cm_drpaddr,
  input  wire  [15:0] gtf_cm_drpdi,
  input  wire   [1:0] gtf_cm_sdm0width,
  input  wire   [1:0] gtf_cm_sdm1width,
  input  wire  [24:0] gtf_cm_sdm0data,
  input  wire  [24:0] gtf_cm_sdm1data,
  input  wire   [2:0] gtf_cm_qpll0refclksel,
  input  wire   [2:0] gtf_cm_qpll1refclksel,
  input  wire   [4:0] gtf_cm_bgrcalovrd,
  input  wire   [4:0] gtf_cm_qpllrsvd2,
  input  wire   [4:0] gtf_cm_qpllrsvd3,
  input  wire   [7:0] gtf_cm_pmarsvd0,
  input  wire   [7:0] gtf_cm_pmarsvd1,
  input  wire   [7:0] gtf_cm_qpll0fbdiv,
  input  wire   [7:0] gtf_cm_qpll1fbdiv,
  input  wire   [7:0] gtf_cm_qpllrsvd1,
  input  wire   [7:0] gtf_cm_qpllrsvd4,
  output wire         gtf_cm_drprdy,
  output wire         gtf_cm_qpll0fbclklost,
  output wire         gtf_cm_qpll0lock,
  output wire         gtf_cm_qpll0outclk,
  output wire         gtf_cm_qpll0outrefclk,
  output wire         gtf_cm_qpll0refclklost,
  output wire         gtf_cm_qpll1fbclklost,
  output wire         gtf_cm_qpll1lock,
  output wire         gtf_cm_qpll1outclk,
  output wire         gtf_cm_qpll1outrefclk,
  output wire         gtf_cm_qpll1refclklost,
  output wire         gtf_cm_refclkoutmonitor0,
  output wire         gtf_cm_refclkoutmonitor1,
  output wire  [14:0] gtf_cm_sdm0testdata,
  output wire  [14:0] gtf_cm_sdm1testdata,
  output wire  [15:0] gtf_cm_drpdo,
  output wire   [1:0] gtf_cm_rxrecclk0sel,
  output wire   [1:0] gtf_cm_rxrecclk1sel,
  output wire   [3:0] gtf_cm_sdm0finalout,
  output wire   [3:0] gtf_cm_sdm1finalout,
  output wire   [7:0] gtf_cm_pmarsvdout0,
  output wire   [7:0] gtf_cm_pmarsvdout1,
  output wire   [7:0] gtf_cm_qplldmonitor0,
  output wire   [7:0] gtf_cm_qplldmonitor1
);


//----{
GTF_COMMON #(
.A_SDM1DATA_HIGH         (A_SDM1DATA_HIGH         ),
.A_SDM1DATA_LOW          (A_SDM1DATA_LOW          ),
.BIAS_CFG0               (BIAS_CFG0               ),
.BIAS_CFG1               (BIAS_CFG1               ),
.BIAS_CFG2               (BIAS_CFG2               ),
.BIAS_CFG3               (BIAS_CFG3               ),
.BIAS_CFG4               (BIAS_CFG4               ),
.BIAS_CFG_RSVD           (BIAS_CFG_RSVD           ),
.COMMON_CFG0             (COMMON_CFG0             ),
.COMMON_CFG1             (COMMON_CFG1             ),
.POR_CFG                 (POR_CFG                 ),
.PPF0_CFG                (PPF0_CFG                ),
.PPF1_CFG                (PPF1_CFG                ),
.QPLL0_CFG0              (QPLL0_CFG0              ),
.QPLL0_CFG1              (QPLL0_CFG1              ),
.QPLL0_CFG1_G3           (QPLL0_CFG1_G3           ),
.QPLL0_CFG2              (QPLL0_CFG2              ),
.QPLL0_CFG2_G3           (QPLL0_CFG2_G3           ),
.QPLL0_CFG3              (QPLL0_CFG3              ),
.QPLL0_CFG4              (QPLL0_CFG4              ),
.QPLL0_CP                (QPLL0_CP                ),
.QPLL0_CP_G3             (QPLL0_CP_G3             ),
.QPLL0_FBDIV             (QPLL0_FBDIV             ),
.QPLL0_FBDIV_G3          (QPLL0_FBDIV_G3          ),
.QPLL0_INIT_CFG0         (QPLL0_INIT_CFG0         ),
.QPLL0_INIT_CFG1         (QPLL0_INIT_CFG1         ),
.QPLL0_LOCK_CFG          (QPLL0_LOCK_CFG          ),
.QPLL0_LOCK_CFG_G3       (QPLL0_LOCK_CFG_G3       ),
.QPLL0_LPF               (QPLL0_LPF               ),
.QPLL0_LPF_G3            (QPLL0_LPF_G3            ),
.QPLL0_REFCLK_DIV        (QPLL0_REFCLK_DIV        ),
.QPLL0_SDM_CFG0          (QPLL0_SDM_CFG0          ),
.QPLL0_SDM_CFG1          (QPLL0_SDM_CFG1          ),
.QPLL0_SDM_CFG2          (QPLL0_SDM_CFG2          ),
.QPLL1_CFG0              (QPLL1_CFG0              ),
.QPLL1_CFG1              (QPLL1_CFG1              ),
.QPLL1_CFG1_G3           (QPLL1_CFG1_G3           ),
.QPLL1_CFG2              (QPLL1_CFG2              ),
.QPLL1_CFG2_G3           (QPLL1_CFG2_G3           ),
.QPLL1_CFG3              (QPLL1_CFG3              ),
.QPLL1_CFG4              (QPLL1_CFG4              ),
.QPLL1_CP                (QPLL1_CP                ),
.QPLL1_CP_G3             (QPLL1_CP_G3             ),
.QPLL1_FBDIV             (QPLL1_FBDIV             ),
.QPLL1_FBDIV_G3          (QPLL1_FBDIV_G3          ),
.QPLL1_INIT_CFG0         (QPLL1_INIT_CFG0         ),
.QPLL1_INIT_CFG1         (QPLL1_INIT_CFG1         ),
.QPLL1_LOCK_CFG          (QPLL1_LOCK_CFG          ),
.QPLL1_LOCK_CFG_G3       (QPLL1_LOCK_CFG_G3       ),
.QPLL1_LPF               (QPLL1_LPF               ),
.QPLL1_LPF_G3            (QPLL1_LPF_G3            ),
.QPLL1_REFCLK_DIV        (QPLL1_REFCLK_DIV        ),
.QPLL1_SDM_CFG0          (QPLL1_SDM_CFG0          ),
.QPLL1_SDM_CFG1          (QPLL1_SDM_CFG1          ),
.QPLL1_SDM_CFG2          (QPLL1_SDM_CFG2          ),
.RSVD_ATTR0              (RSVD_ATTR0              ),
.RSVD_ATTR1              (RSVD_ATTR1              ),
.RSVD_ATTR2              (RSVD_ATTR2              ),
.RSVD_ATTR3              (RSVD_ATTR3              ),
.RXRECCLKOUT0_SEL        (RXRECCLKOUT0_SEL        ),
.RXRECCLKOUT1_SEL        (RXRECCLKOUT1_SEL        ),
.SDM0INITSEED0_0         (SDM0INITSEED0_0         ),
.SDM0INITSEED0_1         (SDM0INITSEED0_1         ),
.SDM1INITSEED0_0         (SDM1INITSEED0_0         ),
.SDM1INITSEED0_1         (SDM1INITSEED0_1         ),
.AEN_QPLL0_FBDIV         (AEN_QPLL0_FBDIV         ),
.AEN_QPLL1_FBDIV         (AEN_QPLL1_FBDIV         ),
.AEN_SDM0TOGGLE          (AEN_SDM0TOGGLE          ),
.AEN_SDM1TOGGLE          (AEN_SDM1TOGGLE          ),
.A_SDM0TOGGLE            (A_SDM0TOGGLE            ),
.A_SDM1TOGGLE            (A_SDM1TOGGLE            ),
.QPLL0CLKOUT_RATE        (QPLL0CLKOUT_RATE        ),
.QPLL0_PCI_EN            (QPLL0_PCI_EN            ),
.QPLL0_RATE_SW_USE_DRP   (QPLL0_RATE_SW_USE_DRP   ),
.QPLL1CLKOUT_RATE        (QPLL1CLKOUT_RATE        ),
.QPLL1_PCI_EN            (QPLL1_PCI_EN            ),
.QPLL1_RATE_SW_USE_DRP   (QPLL1_RATE_SW_USE_DRP   ),
.SARC_ENB                (SARC_ENB                ),
.SARC_SEL                (SARC_SEL                ),
.SIM_MODE                (SIM_MODE                ),
.SIM_RESET_SPEEDUP       (SIM_RESET_SPEEDUP       )
) gtf_common_inst(
.BGBYPASSB          (gtf_cm_bgbypassb          ),
.BGMONITORENB       (gtf_cm_bgmonitorenb       ),
.BGPDB              (gtf_cm_bgpdb              ),
.BGRCALOVRDENB      (gtf_cm_bgrcalovrdenb      ),
.DRPCLK             (gtf_cm_drpclk             ),
.DRPEN              (gtf_cm_drpen              ),
.DRPWE              (gtf_cm_drpwe              ),
.GTGREFCLK0         (gtf_cm_gtgrefclk0         ),
.GTGREFCLK1         (gtf_cm_gtgrefclk1         ),
.GTNORTHREFCLK00    (gtf_cm_gtnorthrefclk00    ),
.GTNORTHREFCLK01    (gtf_cm_gtnorthrefclk01    ),
.GTNORTHREFCLK10    (gtf_cm_gtnorthrefclk10    ),
.GTNORTHREFCLK11    (gtf_cm_gtnorthrefclk11    ),
.GTREFCLK00         (gtf_cm_gtrefclk00         ),
.GTREFCLK01         (gtf_cm_gtrefclk01         ),
.GTREFCLK10         (gtf_cm_gtrefclk10         ),
.GTREFCLK11         (gtf_cm_gtrefclk11         ),
.GTSOUTHREFCLK00    (gtf_cm_gtsouthrefclk00    ),
.GTSOUTHREFCLK01    (gtf_cm_gtsouthrefclk01    ),
.GTSOUTHREFCLK10    (gtf_cm_gtsouthrefclk10    ),
.GTSOUTHREFCLK11    (gtf_cm_gtsouthrefclk11    ),
.QPLL0CLKRSVD0      (gtf_cm_qpll0clkrsvd0      ),
.QPLL0CLKRSVD1      (gtf_cm_qpll0clkrsvd1      ),
.QPLL0LOCKDETCLK    (gtf_cm_qpll0lockdetclk    ),
.QPLL0LOCKEN        (gtf_cm_qpll0locken        ),
.QPLL0PD            (gtf_cm_qpll0pd            ),
.QPLL0RESET         (gtf_cm_qpll0reset         ),
.QPLL1CLKRSVD0      (gtf_cm_qpll1clkrsvd0      ),
.QPLL1CLKRSVD1      (gtf_cm_qpll1clkrsvd1      ),
.QPLL1LOCKDETCLK    (gtf_cm_qpll1lockdetclk    ),
.QPLL1LOCKEN        (gtf_cm_qpll1locken        ),
.QPLL1PD            (gtf_cm_qpll1pd            ),
.QPLL1RESET         (gtf_cm_qpll1reset         ),
.RCALENB            (gtf_cm_rcalenb            ),
.SDM0RESET          (gtf_cm_sdm0reset          ),
.SDM0TOGGLE         (gtf_cm_sdm0toggle         ),
.SDM1RESET          (gtf_cm_sdm1reset          ),
.SDM1TOGGLE         (gtf_cm_sdm1toggle         ),
.DRPADDR            (gtf_cm_drpaddr            ),
.DRPDI              (gtf_cm_drpdi              ),
.SDM0WIDTH          (gtf_cm_sdm0width          ),
.SDM1WIDTH          (gtf_cm_sdm1width          ),
.SDM0DATA           (gtf_cm_sdm0data           ),
.SDM1DATA           (gtf_cm_sdm1data           ),
.QPLL0REFCLKSEL     (gtf_cm_qpll0refclksel     ),
.QPLL1REFCLKSEL     (gtf_cm_qpll1refclksel     ),
.BGRCALOVRD         (gtf_cm_bgrcalovrd         ),
.QPLLRSVD2          (gtf_cm_qpllrsvd2          ),
.QPLLRSVD3          (gtf_cm_qpllrsvd3          ),
.PMARSVD0           (gtf_cm_pmarsvd0           ),
.PMARSVD1           (gtf_cm_pmarsvd1           ),
.QPLL0FBDIV         (gtf_cm_qpll0fbdiv         ),
.QPLL1FBDIV         (gtf_cm_qpll1fbdiv         ),
.QPLLRSVD1          (gtf_cm_qpllrsvd1          ),
.QPLLRSVD4          (gtf_cm_qpllrsvd4          ),
.DRPRDY             (gtf_cm_drprdy             ),
.QPLL0FBCLKLOST     (gtf_cm_qpll0fbclklost     ),
.QPLL0LOCK          (gtf_cm_qpll0lock          ),
.QPLL0OUTCLK        (gtf_cm_qpll0outclk        ),
.QPLL0OUTREFCLK     (gtf_cm_qpll0outrefclk     ),
.QPLL0REFCLKLOST    (gtf_cm_qpll0refclklost    ),
.QPLL1FBCLKLOST     (gtf_cm_qpll1fbclklost     ),
.QPLL1LOCK          (gtf_cm_qpll1lock          ),
.QPLL1OUTCLK        (gtf_cm_qpll1outclk        ),
.QPLL1OUTREFCLK     (gtf_cm_qpll1outrefclk     ),
.QPLL1REFCLKLOST    (gtf_cm_qpll1refclklost    ),
.REFCLKOUTMONITOR0  (gtf_cm_refclkoutmonitor0  ),
.REFCLKOUTMONITOR1  (gtf_cm_refclkoutmonitor1  ),
.SDM0TESTDATA       (gtf_cm_sdm0testdata       ),
.SDM1TESTDATA       (gtf_cm_sdm1testdata       ),
.DRPDO              (gtf_cm_drpdo              ),
.RXRECCLK0SEL       (gtf_cm_rxrecclk0sel       ),
.RXRECCLK1SEL       (gtf_cm_rxrecclk1sel       ),
.SDM0FINALOUT       (gtf_cm_sdm0finalout       ),
.SDM1FINALOUT       (gtf_cm_sdm1finalout       ),
.PMARSVDOUT0        (gtf_cm_pmarsvdout0        ),
.PMARSVDOUT1        (gtf_cm_pmarsvdout1        ),
.QPLLDMONITOR0      (gtf_cm_qplldmonitor0      ),
.QPLLDMONITOR1      (gtf_cm_qplldmonitor1      )
);
//----}


endmodule
`default_nettype wire
//------}
