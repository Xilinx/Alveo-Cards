/*
Copyright (c) 2023, Advanced Micro Devices, Inc. All rights reserved.
SPDX-License-Identifier: MIT
*/

//------------------------------------------------------------------------------


//------{
`timescale 1fs/1fs
`default_nettype none
(* DowngradeIPIdentifiedWarnings="yes" *)
module gtfwizard_0 (
  input  wire       gtwiz_reset_clk_freerun_in,
  input  wire       gtwiz_reset_all_in,
  input  wire       gtwiz_reset_tx_pll_and_datapath_in,
  input  wire       gtwiz_reset_tx_datapath_in,
  input  wire       gtwiz_reset_rx_pll_and_datapath_in,
  input  wire       gtwiz_reset_rx_datapath_in,
  output wire       gtwiz_reset_rx_cdr_stable_out,
  output wire       gtwiz_reset_tx_done_out,
  output wire       gtwiz_reset_rx_done_out,
  output wire       gtwiz_pllreset_rx_out,
  output wire       gtwiz_pllreset_tx_out,
  input  wire       plllock_tx_in,
  input  wire       plllock_rx_in,
  input  wire       gtf_ch_cdrstepdir,
  input  wire       gtf_ch_cdrstepsq,
  input  wire       gtf_ch_cdrstepsx,
  input  wire       gtf_ch_cfgreset,
  input  wire       gtf_ch_clkrsvd0,
  input  wire       gtf_ch_clkrsvd1,
  input  wire       gtf_ch_cpllfreqlock,
  input  wire       gtf_ch_cplllockdetclk,
  input  wire       gtf_ch_cplllocken,
  input  wire       gtf_ch_cpllpd,
  input  wire       gtf_ch_cpllreset,
  input  wire       gtf_ch_ctltxresendpause,
  input  wire       gtf_ch_dmonfiforeset,
  input  wire       gtf_ch_dmonitorclk,
  input  wire       gtf_ch_drpclk,
  input  wire       gtf_ch_drprst,
  input  wire       gtf_ch_eyescanreset,
  input  wire       gtf_ch_eyescantrigger,
  input  wire       gtf_ch_freqos,
  input  wire       gtf_ch_gtfrxn,
  input  wire       gtf_ch_gtfrxp,
  input  wire       gtf_ch_gtgrefclk,
  input  wire       gtf_ch_gtnorthrefclk0,
  input  wire       gtf_ch_gtnorthrefclk1,
  input  wire       gtf_ch_gtrefclk0,
  input  wire       gtf_ch_gtrefclk1,
  input  wire       gtf_ch_gtrxresetsel,
  input  wire       gtf_ch_gtsouthrefclk0,
  input  wire       gtf_ch_gtsouthrefclk1,
  input  wire       gtf_ch_gttxresetsel,
  input  wire       gtf_ch_incpctrl,
  input  wire       gtf_ch_qpll0clk,
  input  wire       gtf_ch_qpll0freqlock,
  input  wire       gtf_ch_qpll0refclk,
  input  wire       gtf_ch_qpll1clk,
  input  wire       gtf_ch_qpll1freqlock,
  input  wire       gtf_ch_qpll1refclk,
  input  wire       gtf_ch_resetovrd,
  input  wire       gtf_ch_rxafecfoken,
  input  wire       gtf_ch_rxcdrfreqreset,
  input  wire       gtf_ch_rxcdrhold,
  input  wire       gtf_ch_rxcdrovrden,
  input  wire       gtf_ch_rxcdrreset,
  input  wire       gtf_ch_rxckcalreset,
  input  wire       gtf_ch_rxdfeagchold,
  input  wire       gtf_ch_rxdfeagcovrden,
  input  wire       gtf_ch_rxdfecfokfen,
  input  wire       gtf_ch_rxdfecfokfpulse,
  input  wire       gtf_ch_rxdfecfokhold,
  input  wire       gtf_ch_rxdfecfokovren,
  input  wire       gtf_ch_rxdfekhhold,
  input  wire       gtf_ch_rxdfekhovrden,
  input  wire       gtf_ch_rxdfelfhold,
  input  wire       gtf_ch_rxdfelfovrden,
  input  wire       gtf_ch_rxdfelpmreset,
  input  wire       gtf_ch_rxdfetap10hold,
  input  wire       gtf_ch_rxdfetap10ovrden,
  input  wire       gtf_ch_rxdfetap11hold,
  input  wire       gtf_ch_rxdfetap11ovrden,
  input  wire       gtf_ch_rxdfetap12hold,
  input  wire       gtf_ch_rxdfetap12ovrden,
  input  wire       gtf_ch_rxdfetap13hold,
  input  wire       gtf_ch_rxdfetap13ovrden,
  input  wire       gtf_ch_rxdfetap14hold,
  input  wire       gtf_ch_rxdfetap14ovrden,
  input  wire       gtf_ch_rxdfetap15hold,
  input  wire       gtf_ch_rxdfetap15ovrden,
  input  wire       gtf_ch_rxdfetap2hold,
  input  wire       gtf_ch_rxdfetap2ovrden,
  input  wire       gtf_ch_rxdfetap3hold,
  input  wire       gtf_ch_rxdfetap3ovrden,
  input  wire       gtf_ch_rxdfetap4hold,
  input  wire       gtf_ch_rxdfetap4ovrden,
  input  wire       gtf_ch_rxdfetap5hold,
  input  wire       gtf_ch_rxdfetap5ovrden,
  input  wire       gtf_ch_rxdfetap6hold,
  input  wire       gtf_ch_rxdfetap6ovrden,
  input  wire       gtf_ch_rxdfetap7hold,
  input  wire       gtf_ch_rxdfetap7ovrden,
  input  wire       gtf_ch_rxdfetap8hold,
  input  wire       gtf_ch_rxdfetap8ovrden,
  input  wire       gtf_ch_rxdfetap9hold,
  input  wire       gtf_ch_rxdfetap9ovrden,
  input  wire       gtf_ch_rxdfeuthold,
  input  wire       gtf_ch_rxdfeutovrden,
  input  wire       gtf_ch_rxdfevphold,
  input  wire       gtf_ch_rxdfevpovrden,
  input  wire       gtf_ch_rxdfexyden,
  input  wire       gtf_ch_rxlpmen,
  input  wire       gtf_ch_rxlpmgchold,
  input  wire       gtf_ch_rxlpmgcovrden,
  input  wire       gtf_ch_rxlpmhfhold,
  input  wire       gtf_ch_rxlpmhfovrden,
  input  wire       gtf_ch_rxlpmlfhold,
  input  wire       gtf_ch_rxlpmlfklovrden,
  input  wire       gtf_ch_rxlpmoshold,
  input  wire       gtf_ch_rxlpmosovrden,
  input  wire       gtf_ch_rxoscalreset,
  input  wire       gtf_ch_rxoshold,
  input  wire       gtf_ch_rxosovrden,
  input  wire       gtf_ch_rxpcsreset,
  input  wire       gtf_ch_rxpmareset,
  input  wire       gtf_ch_rxpolarity,
  input  wire       gtf_ch_rxprbscntreset,
  input  wire       gtf_ch_rxslipoutclk,
  input  wire   gtf_ch_rxslippma,
  input  wire       gtf_ch_rxtermination,
  input  wire       gtf_ch_rxuserrdy,
  input  wire       gtf_ch_txaxisterr,
  input  wire       gtf_ch_txaxistpoison,
  input  wire       gtf_ch_txaxistvalid,
  input  wire       gtf_ch_txdccforcestart,
  input  wire       gtf_ch_txdccreset,
  input  wire       gtf_ch_txelecidle,
  input  wire       gtf_ch_txgbseqsync,
  input  wire       gtf_ch_txmuxdcdexhold,
  input  wire       gtf_ch_txmuxdcdorwren,
  input  wire       gtf_ch_txpcsreset,
  input  wire       gtf_ch_txpippmen,
  input  wire       gtf_ch_txpippmovrden,
  input  wire       gtf_ch_txpippmpd,
  input  wire       gtf_ch_txpippmsel,
  input  wire       gtf_ch_txpisopd,
  input  wire       gtf_ch_txpmareset,
  input  wire       gtf_ch_txpolarity,
  input  wire       gtf_ch_txprbsforceerr,
  input  wire       gtf_ch_txuserrdy,
  input  wire [15:0]      gtf_ch_gtrsvd,
  input  wire [15:0]      gtf_ch_pcsrsvdin,
  input  wire [19:0]      gtf_ch_tstin,
  input  wire [1:0]       gtf_ch_rxelecidlemode,
  input  wire [1:0]       gtf_ch_rxmonitorsel,
  input  wire [1:0]       gtf_ch_rxpd,
  input  wire [1:0]       gtf_ch_rxpllclksel,
  input  wire [1:0]       gtf_ch_rxsysclksel,
  input  wire [1:0]       gtf_ch_txaxistsof,
  input  wire [1:0]       gtf_ch_txpd,
  input  wire [1:0]       gtf_ch_txpllclksel,
  input  wire [1:0]       gtf_ch_txsysclksel,
  input  wire [2:0]       gtf_ch_cpllrefclksel,
  input  wire [2:0]       gtf_ch_rxoutclksel,
  input  wire [2:0]       gtf_ch_txoutclksel,
  input  wire [39:0]      gtf_ch_txrawdata,
  input  wire [3:0]       gtf_ch_rxdfecfokfcnum,
  input  wire [3:0]       gtf_ch_rxprbssel,
  input  wire [3:0]       gtf_ch_txprbssel,
  input  wire [4:0]       gtf_ch_txaxistterm,
  input  wire [4:0]       gtf_ch_txdiffctrl,
  input  wire [4:0]       gtf_ch_txpippmstepsize,
  input  wire [4:0]       gtf_ch_txpostcursor,
  input  wire [4:0]       gtf_ch_txprecursor,
  input  wire [63:0]      gtf_ch_txaxistdata,
  input  wire [6:0]       gtf_ch_rxckcalstart,
  input  wire [6:0]       gtf_ch_txmaincursor,
  input  wire [7:0]       gtf_ch_txaxistlast,
  input  wire [7:0]       gtf_ch_txaxistpre,
  input  wire [8:0]       gtf_ch_ctlrxpauseack,
  input  wire [8:0]       gtf_ch_ctltxpausereq,
  output wire       gtf_ch_cpllfbclklost,
  output wire       gtf_ch_cplllock,
  output wire       gtf_ch_cpllrefclklost,
  output wire       gtf_ch_dmonitoroutclk,
  output wire       gtf_ch_eyescandataerror,
  output wire       gtf_ch_gtftxn,
  output wire       gtf_ch_gtftxp,
  output wire       gtf_ch_gtpowergood,
  output wire       gtf_ch_gtrefclkmonitor,
  output wire       gtf_ch_resetexception,
  output wire       gtf_ch_rxaxisterr,
  output wire       gtf_ch_rxaxistvalid,
  output wire       gtf_ch_rxbitslip,
  output wire       gtf_ch_rxcdrlock,
  output wire       gtf_ch_rxcdrphdone,
  output wire       gtf_ch_rxckcaldone,
  output wire       gtf_ch_rxelecidle,
  output wire       gtf_ch_rxgbseqstart,
  output wire       gtf_ch_rxosintdone,
  output wire       gtf_ch_rxosintstarted,
  output wire       gtf_ch_rxosintstrobedone,
  output wire       gtf_ch_rxosintstrobestarted,
  output wire       gtf_ch_rxoutclk,
  output wire       gtf_ch_rxoutclkfabric,
  output wire       gtf_ch_rxoutclkpcs,
  output wire       gtf_ch_rxphalignerr,
  output wire       gtf_ch_rxpmaresetdone,
  output wire       gtf_ch_rxprbserr,
  output wire       gtf_ch_rxprbslocked,
  output wire       gtf_ch_rxprgdivresetdone,
  output wire       gtf_ch_rxptpsop,
  output wire       gtf_ch_rxptpsoppos,
  output wire       gtf_ch_rxrecclkout,
  output wire       gtf_ch_rxresetdone,
  output wire       gtf_ch_rxslipdone,
  output wire       gtf_ch_rxslipoutclkrdy,
  output wire       gtf_ch_rxslippmardy,
  output wire       gtf_ch_rxsyncdone,




  output wire       gtf_ch_statrxblocklock,

  output wire       gtf_ch_statrxfcserr,

  input  wire       gtf_ch_ctltxsendlfi,
  input  wire       gtf_ch_ctltxsendrfi,
  input  wire       gtf_ch_ctltxsendidle,


  output wire       gtf_ch_statrxhiber,
  output wire       gtf_ch_statrxstatus,
  output wire       gtf_ch_statrxpkterr,
  output wire       gtf_ch_statrxbadpreamble,
  output wire       gtf_ch_statrxbadsfd,
  output wire       gtf_ch_statrxgotsignalos,
  output wire       gtf_ch_statrxbadcode,
  output wire       gtf_ch_statrxstompedfcs,
  output wire       gtf_ch_statrxframingerr,
  output wire       gtf_ch_statrxtruncated,
  output wire [3:0]      gtf_ch_statrxbytes,
  output wire       gtf_ch_statrxpkt,
  output wire       gtf_ch_statrxbadfcs,
  output wire       gtf_ch_statrxunicast,
  output wire       gtf_ch_statrxbroadcast,
  output wire       gtf_ch_statrxvlan,
  output wire   gtf_ch_statrxinrangeerr,
  output wire [8:0]  gtf_ch_statrxpausevalid,
  output wire [8:0]  gtf_ch_statrxpausereq,
  output wire [8:0]  gtf_ch_statrxpausequanta,
  output wire [3:0]  gtf_ch_stattxbytes,
  output wire        gtf_ch_stattxpkt,
  output wire        gtf_ch_stattxpkterr,
  output wire        gtf_ch_stattxbadfcs,
  output wire        gtf_ch_stattxunicast,
  output wire        gtf_ch_stattxbroadcast,
  output wire        gtf_ch_stattxmulticast,
  output wire        gtf_ch_stattxvlan,
  output wire        gtf_ch_statrxmulticast,
  input  wire [2:0]  gtf_ch_loopback,
  output wire       gtf_ch_statrxinternallocalfault,
  output wire       gtf_ch_statrxlocalfault,


  output wire       gtf_ch_statrxreceivedlocalfault,
  output wire       gtf_ch_statrxremotefault,


  output wire       gtf_ch_statrxtestpatternmismatch,


  output wire       gtf_ch_statrxvalidctrlcode,

  output wire       gtf_ch_stattxfcserr,
  output wire       gtf_ch_txaxistready,
  output wire       gtf_ch_txdccdone,
  output wire       gtf_ch_txgbseqstart,
  output wire       gtf_ch_txoutclk,
  output wire       gtf_ch_txoutclkfabric,
  output wire       gtf_ch_txoutclkpcs,
  output wire       gtf_ch_txpmaresetdone,
  output wire       gtf_ch_txprgdivresetdone,
  output wire       gtf_ch_txptpsop,
  output wire       gtf_ch_txptpsoppos,
  output wire       gtf_ch_txresetdone,
  output wire       gtf_ch_txsyncdone,
  output wire            gtf_ch_txaxistcanstart,
  output wire            gtf_ch_rxinvalidstart,
  output wire            gtf_ch_txunfout,
  output wire     gtwiz_buffbypass_rx_done_out,
  output wire [15:0]     gtf_ch_pcsrsvdout,
  output wire [15:0]     gtf_ch_pinrsrvdas,
  output wire [1:0]      gtf_ch_rxaxistsof,
  output wire [39:0]     gtf_ch_rxrawdata,

  output wire [4:0]      gtf_ch_rxaxistterm,
  output wire [63:0]     gtf_ch_rxaxistdata,
  output wire [7:0]      gtf_ch_rxaxistlast,
  output wire [7:0]      gtf_ch_rxaxistpre,
  output wire [7:0]      gtf_ch_rxmonitorout,
  output wire [8:0]      gtf_ch_stattxpausevalid,
  output wire       gtf_ch_gttxreset_out,
  output wire       gtwiz_buffbypass_tx_done_out,
  output wire       gtf_txusrclk2_out,
  output wire       gtf_rxusrclk2_out
);

//------{
`ifdef XIL_TIMING
  parameter LOC = "UNPLACED";
`endif

`include "gtfwizard_0_rules_output.vh" 
//------}



gtfwizard_0_top # (
.ACJTAG_DEBUG_MODE               (ACJTAG_DEBUG_MODE               ),
.ACJTAG_MODE                     (ACJTAG_MODE                     ),
.ACJTAG_RESET                    (ACJTAG_RESET                    ),
.ADAPT_CFG0                      (ADAPT_CFG0                      ),
.ADAPT_CFG1                      (ADAPT_CFG1                      ),
.ADAPT_CFG2                      (ADAPT_CFG2                      ),
.AEN_QPLL0_FBDIV                 (AEN_QPLL0_FBDIV                 ),
.AEN_QPLL1_FBDIV                 (AEN_QPLL1_FBDIV                 ),
.AEN_SDM0TOGGLE                  (AEN_SDM0TOGGLE                  ),
.AEN_SDM1TOGGLE                  (AEN_SDM1TOGGLE                  ),
.A_RXOSCALRESET                  (A_RXOSCALRESET                  ),
.A_RXPROGDIVRESET                (A_RXPROGDIVRESET                ),
.A_RXTERMINATION                 (A_RXTERMINATION                 ),
.A_SDM0TOGGLE                    (A_SDM0TOGGLE                    ),
.A_SDM1DATA_HIGH                 (A_SDM1DATA_HIGH                 ),
.A_SDM1DATA_LOW                  (A_SDM1DATA_LOW                  ),
.A_SDM1TOGGLE                    (A_SDM1TOGGLE                    ),
.A_TXDIFFCTRL                    (A_TXDIFFCTRL                    ),
.A_TXPROGDIVRESET                (A_TXPROGDIVRESET                ),
.BIAS_CFG0                       (BIAS_CFG0                       ),
.BIAS_CFG1                       (BIAS_CFG1                       ),
.BIAS_CFG2                       (BIAS_CFG2                       ),
.BIAS_CFG3                       (BIAS_CFG3                       ),
.BIAS_CFG4                       (BIAS_CFG4                       ),
.BIAS_CFG_RSVD                   (BIAS_CFG_RSVD                   ),
.CBCC_DATA_SOURCE_SEL            (CBCC_DATA_SOURCE_SEL            ),
.CDR_SWAP_MODE_EN                (CDR_SWAP_MODE_EN                ),
.CFOK_PWRSVE_EN                  (CFOK_PWRSVE_EN                  ),
.CH_HSPMUX                       (CH_HSPMUX                       ),
.CKCAL1_CFG_0                    (CKCAL1_CFG_0                    ),
.CKCAL1_CFG_1                    (CKCAL1_CFG_1                    ),
.CKCAL1_CFG_2                    (CKCAL1_CFG_2                    ),
.CKCAL1_CFG_3                    (CKCAL1_CFG_3                    ),
.CKCAL2_CFG_0                    (CKCAL2_CFG_0                    ),
.CKCAL2_CFG_1                    (CKCAL2_CFG_1                    ),
.CKCAL2_CFG_2                    (CKCAL2_CFG_2                    ),
.CKCAL2_CFG_3                    (CKCAL2_CFG_3                    ),
.CKCAL2_CFG_4                    (CKCAL2_CFG_4                    ),
.COMMON_CFG0                     (COMMON_CFG0                     ),
.COMMON_CFG1                     (COMMON_CFG1                     ),
.CPLL_CFG0                       (CPLL_CFG0                       ),
.CPLL_CFG1                       (CPLL_CFG1                       ),
.CPLL_CFG2                       (CPLL_CFG2                       ),
.CPLL_CFG3                       (CPLL_CFG3                       ),
.CPLL_FBDIV                      (CPLL_FBDIV                      ),
.CPLL_FBDIV_45                   (CPLL_FBDIV_45                   ),
.CPLL_INIT_CFG0                  (CPLL_INIT_CFG0                  ),
.CPLL_LOCK_CFG                   (CPLL_LOCK_CFG                   ),
.CPLL_REFCLK_DIV                 (CPLL_REFCLK_DIV                 ),
.CTLE3_OCAP_EXT_CTRL             (CTLE3_OCAP_EXT_CTRL             ),
.CTLE3_OCAP_EXT_EN               (CTLE3_OCAP_EXT_EN               ),
.DDI_CTRL                        (DDI_CTRL                        ),
.DDI_REALIGN_WAIT                (DDI_REALIGN_WAIT                ),
.DELAY_ELEC                      (DELAY_ELEC                      ),
.DMONITOR_CFG0                   (DMONITOR_CFG0                   ),
.DMONITOR_CFG1                   (DMONITOR_CFG1                   ),
.ES_CLK_PHASE_SEL                (ES_CLK_PHASE_SEL                ),
.ES_CONTROL                      (ES_CONTROL                      ),
.ES_ERRDET_EN                    (ES_ERRDET_EN                    ),
.ES_EYE_SCAN_EN                  (ES_EYE_SCAN_EN                  ),
.ES_HORZ_OFFSET                  (ES_HORZ_OFFSET                  ),
.ES_PRESCALE                     (ES_PRESCALE                     ),
.ES_QUALIFIER0                   (ES_QUALIFIER0                   ),
.ES_QUALIFIER1                   (ES_QUALIFIER1                   ),
.ES_QUALIFIER2                   (ES_QUALIFIER2                   ),
.ES_QUALIFIER3                   (ES_QUALIFIER3                   ),
.ES_QUALIFIER4                   (ES_QUALIFIER4                   ),
.ES_QUALIFIER5                   (ES_QUALIFIER5                   ),
.ES_QUALIFIER6                   (ES_QUALIFIER6                   ),
.ES_QUALIFIER7                   (ES_QUALIFIER7                   ),
.ES_QUALIFIER8                   (ES_QUALIFIER8                   ),
.ES_QUALIFIER9                   (ES_QUALIFIER9                   ),
.ES_QUAL_MASK0                   (ES_QUAL_MASK0                   ),
.ES_QUAL_MASK1                   (ES_QUAL_MASK1                   ),
.ES_QUAL_MASK2                   (ES_QUAL_MASK2                   ),
.ES_QUAL_MASK3                   (ES_QUAL_MASK3                   ),
.ES_QUAL_MASK4                   (ES_QUAL_MASK4                   ),
.ES_QUAL_MASK5                   (ES_QUAL_MASK5                   ),
.ES_QUAL_MASK6                   (ES_QUAL_MASK6                   ),
.ES_QUAL_MASK7                   (ES_QUAL_MASK7                   ),
.ES_QUAL_MASK8                   (ES_QUAL_MASK8                   ),
.ES_QUAL_MASK9                   (ES_QUAL_MASK9                   ),
.ES_SDATA_MASK0                  (ES_SDATA_MASK0                  ),
.ES_SDATA_MASK1                  (ES_SDATA_MASK1                  ),
.ES_SDATA_MASK2                  (ES_SDATA_MASK2                  ),
.ES_SDATA_MASK3                  (ES_SDATA_MASK3                  ),
.ES_SDATA_MASK4                  (ES_SDATA_MASK4                  ),
.ES_SDATA_MASK5                  (ES_SDATA_MASK5                  ),
.ES_SDATA_MASK6                  (ES_SDATA_MASK6                  ),
.ES_SDATA_MASK7                  (ES_SDATA_MASK7                  ),
.ES_SDATA_MASK8                  (ES_SDATA_MASK8                  ),
.ES_SDATA_MASK9                  (ES_SDATA_MASK9                  ),
.EYESCAN_VP_RANGE                (EYESCAN_VP_RANGE                ),
.EYE_SCAN_SWAP_EN                (EYE_SCAN_SWAP_EN                ),
.FTS_DESKEW_SEQ_ENABLE           (FTS_DESKEW_SEQ_ENABLE           ),
.FTS_LANE_DESKEW_CFG             (FTS_LANE_DESKEW_CFG             ),
.FTS_LANE_DESKEW_EN              (FTS_LANE_DESKEW_EN              ),
.GEARBOX_MODE                    (GEARBOX_MODE                    ),
.ISCAN_CK_PH_SEL2                (ISCAN_CK_PH_SEL2                ),
.LOCAL_MASTER                    (LOCAL_MASTER                    ),
.LPBK_BIAS_CTRL                  (LPBK_BIAS_CTRL                  ),
.LPBK_EN_RCAL_B                  (LPBK_EN_RCAL_B                  ),
.LPBK_EXT_RCAL                   (LPBK_EXT_RCAL                   ),
.LPBK_IND_CTRL0                  (LPBK_IND_CTRL0                  ),
.LPBK_IND_CTRL1                  (LPBK_IND_CTRL1                  ),
.LPBK_IND_CTRL2                  (LPBK_IND_CTRL2                  ),
.LPBK_RG_CTRL                    (LPBK_RG_CTRL                    ),
.MAC_CFG0                        (MAC_CFG0                        ),
.MAC_CFG1                        (MAC_CFG1                        ),
.MAC_CFG10                       (MAC_CFG10                       ),
.MAC_CFG11                       (MAC_CFG11                       ),
.MAC_CFG12                       (MAC_CFG12                       ),
.MAC_CFG13                       (MAC_CFG13                       ),
.MAC_CFG14                       (MAC_CFG14                       ),
.MAC_CFG15                       (MAC_CFG15                       ),
.MAC_CFG2                        (MAC_CFG2                        ),
.MAC_CFG3                        (MAC_CFG3                        ),
.MAC_CFG4                        (MAC_CFG4                        ),
.MAC_CFG5                        (MAC_CFG5                        ),
.MAC_CFG6                        (MAC_CFG6                        ),
.MAC_CFG7                        (MAC_CFG7                        ),
.MAC_CFG8                        (MAC_CFG8                        ),
.MAC_CFG9                        (MAC_CFG9                        ),
.PCS_RSVD0                       (PCS_RSVD0                       ),
.PD_TRANS_TIME_FROM_P2           (PD_TRANS_TIME_FROM_P2           ),
.PD_TRANS_TIME_NONE_P2           (PD_TRANS_TIME_NONE_P2           ),
.PD_TRANS_TIME_TO_P2             (PD_TRANS_TIME_TO_P2             ),
.POR_CFG                         (POR_CFG                         ),
.PPF0_CFG                        (PPF0_CFG                        ),
.PPF1_CFG                        (PPF1_CFG                        ),
.PREIQ_FREQ_BST                  (PREIQ_FREQ_BST                  ),
.QPLL0CLKOUT_RATE                (QPLL0CLKOUT_RATE                ),
.QPLL0_CFG0                      (QPLL0_CFG0                      ),
.QPLL0_CFG1                      (QPLL0_CFG1                      ),
.QPLL0_CFG1_G3                   (QPLL0_CFG1_G3                   ),
.QPLL0_CFG2                      (QPLL0_CFG2                      ),
.QPLL0_CFG2_G3                   (QPLL0_CFG2_G3                   ),
.QPLL0_CFG3                      (QPLL0_CFG3                      ),
.QPLL0_CFG4                      (QPLL0_CFG4                      ),
.QPLL0_CP                        (QPLL0_CP                        ),
.QPLL0_CP_G3                     (QPLL0_CP_G3                     ),
.QPLL0_FBDIV                     (QPLL0_FBDIV                     ),
.QPLL0_FBDIV_G3                  (QPLL0_FBDIV_G3                  ),
.QPLL0_INIT_CFG0                 (QPLL0_INIT_CFG0                 ),
.QPLL0_INIT_CFG1                 (QPLL0_INIT_CFG1                 ),
.QPLL0_LOCK_CFG                  (QPLL0_LOCK_CFG                  ),
.QPLL0_LOCK_CFG_G3               (QPLL0_LOCK_CFG_G3               ),
.QPLL0_LPF                       (QPLL0_LPF                       ),
.QPLL0_LPF_G3                    (QPLL0_LPF_G3                    ),
.QPLL0_PCI_EN                    (QPLL0_PCI_EN                    ),
.QPLL0_RATE_SW_USE_DRP           (QPLL0_RATE_SW_USE_DRP           ),
.QPLL0_REFCLK_DIV                (QPLL0_REFCLK_DIV                ),
.QPLL0_SDM_CFG0                  (QPLL0_SDM_CFG0                  ),
.QPLL0_SDM_CFG1                  (QPLL0_SDM_CFG1                  ),
.QPLL0_SDM_CFG2                  (QPLL0_SDM_CFG2                  ),
.QPLL1CLKOUT_RATE                (QPLL1CLKOUT_RATE                ),
.QPLL1_CFG0                      (QPLL1_CFG0                      ),
.QPLL1_CFG1                      (QPLL1_CFG1                      ),
.QPLL1_CFG1_G3                   (QPLL1_CFG1_G3                   ),
.QPLL1_CFG2                      (QPLL1_CFG2                      ),
.QPLL1_CFG2_G3                   (QPLL1_CFG2_G3                   ),
.QPLL1_CFG3                      (QPLL1_CFG3                      ),
.QPLL1_CFG4                      (QPLL1_CFG4                      ),
.QPLL1_CP                        (QPLL1_CP                        ),
.QPLL1_CP_G3                     (QPLL1_CP_G3                     ),
.QPLL1_FBDIV                     (QPLL1_FBDIV                     ),
.QPLL1_FBDIV_G3                  (QPLL1_FBDIV_G3                  ),
.QPLL1_INIT_CFG0                 (QPLL1_INIT_CFG0                 ),
.QPLL1_INIT_CFG1                 (QPLL1_INIT_CFG1                 ),
.QPLL1_LOCK_CFG                  (QPLL1_LOCK_CFG                  ),
.QPLL1_LOCK_CFG_G3               (QPLL1_LOCK_CFG_G3               ),
.QPLL1_LPF                       (QPLL1_LPF                       ),
.QPLL1_LPF_G3                    (QPLL1_LPF_G3                    ),
.QPLL1_PCI_EN                    (QPLL1_PCI_EN                    ),
.QPLL1_RATE_SW_USE_DRP           (QPLL1_RATE_SW_USE_DRP           ),
.QPLL1_REFCLK_DIV                (QPLL1_REFCLK_DIV                ),
.QPLL1_SDM_CFG0                  (QPLL1_SDM_CFG0                  ),
.QPLL1_SDM_CFG1                  (QPLL1_SDM_CFG1                  ),
.QPLL1_SDM_CFG2                  (QPLL1_SDM_CFG2                  ),
.RAW_MAC_CFG                     (RAW_MAC_CFG                     ),
.RCLK_SIPO_DLY_ENB               (RCLK_SIPO_DLY_ENB               ),
.RCLK_SIPO_INV_EN                (RCLK_SIPO_INV_EN                ),
.RCO_NEW_MAC_CFG0                (RCO_NEW_MAC_CFG0                ),
.RCO_NEW_MAC_CFG1                (RCO_NEW_MAC_CFG1                ),
.RCO_NEW_MAC_CFG2                (RCO_NEW_MAC_CFG2                ),
.RCO_NEW_MAC_CFG3                (RCO_NEW_MAC_CFG3                ),
.RCO_NEW_RAW_CFG0                (RCO_NEW_RAW_CFG0                ),
.RCO_NEW_RAW_CFG1                (RCO_NEW_RAW_CFG1                ),
.RCO_NEW_RAW_CFG2                (RCO_NEW_RAW_CFG2                ),
.RCO_NEW_RAW_CFG3                (RCO_NEW_RAW_CFG3                ),
.RSVD_ATTR0                      (RSVD_ATTR0                      ),
.RSVD_ATTR1                      (RSVD_ATTR1                      ),
.RSVD_ATTR2                      (RSVD_ATTR2                      ),
.RSVD_ATTR3                      (RSVD_ATTR3                      ),
.RTX_BUF_CML_CTRL                (RTX_BUF_CML_CTRL                ),
.RTX_BUF_TERM_CTRL               (RTX_BUF_TERM_CTRL               ),
.RXBUFRESET_TIME                 (RXBUFRESET_TIME                 ),
.RXBUF_EN                        (RXBUF_EN                        ),
.RXCDRFREQRESET_TIME             (RXCDRFREQRESET_TIME             ),
.RXCDRPHRESET_TIME               (RXCDRPHRESET_TIME               ),
.RXCDR_CFG0                      (RXCDR_CFG0                      ),
.RXCDR_CFG1                      (RXCDR_CFG1                      ),
.RXCDR_CFG2                      (RXCDR_CFG2                      ),
.RXCDR_CFG3                      (RXCDR_CFG3                      ),
.RXCDR_CFG4                      (RXCDR_CFG4                      ),
.RXCDR_CFG5                      (RXCDR_CFG5                      ),
.RXCDR_FR_RESET_ON_EIDLE         (RXCDR_FR_RESET_ON_EIDLE         ),
.RXCDR_HOLD_DURING_EIDLE         (RXCDR_HOLD_DURING_EIDLE         ),
.RXCDR_LOCK_CFG0                 (RXCDR_LOCK_CFG0                 ),
.RXCDR_LOCK_CFG1                 (RXCDR_LOCK_CFG1                 ),
.RXCDR_LOCK_CFG2                 (RXCDR_LOCK_CFG2                 ),
.RXCDR_LOCK_CFG3                 (RXCDR_LOCK_CFG3                 ),
.RXCDR_LOCK_CFG4                 (RXCDR_LOCK_CFG4                 ),
.RXCDR_PH_RESET_ON_EIDLE         (RXCDR_PH_RESET_ON_EIDLE         ),
.RXCFOK_CFG0                     (RXCFOK_CFG0                     ),
.RXCFOK_CFG1                     (RXCFOK_CFG1                     ),
.RXCFOK_CFG2                     (RXCFOK_CFG2                     ),
.RXCKCAL1_IQ_LOOP_RST_CFG        (RXCKCAL1_IQ_LOOP_RST_CFG        ),
.RXCKCAL1_I_LOOP_RST_CFG         (RXCKCAL1_I_LOOP_RST_CFG         ),
.RXCKCAL1_Q_LOOP_RST_CFG         (RXCKCAL1_Q_LOOP_RST_CFG         ),
.RXCKCAL2_DX_LOOP_RST_CFG        (RXCKCAL2_DX_LOOP_RST_CFG        ),
.RXCKCAL2_D_LOOP_RST_CFG         (RXCKCAL2_D_LOOP_RST_CFG         ),
.RXCKCAL2_S_LOOP_RST_CFG         (RXCKCAL2_S_LOOP_RST_CFG         ),
.RXCKCAL2_X_LOOP_RST_CFG         (RXCKCAL2_X_LOOP_RST_CFG         ),
.RXDFELPMRESET_TIME              (RXDFELPMRESET_TIME              ),
.RXDFELPM_KL_CFG0                (RXDFELPM_KL_CFG0                ),
.RXDFELPM_KL_CFG1                (RXDFELPM_KL_CFG1                ),
.RXDFELPM_KL_CFG2                (RXDFELPM_KL_CFG2                ),
.RXDFE_CFG0                      (RXDFE_CFG0                      ),
.RXDFE_CFG1                      (RXDFE_CFG1                      ),
.RXDFE_GC_CFG0                   (RXDFE_GC_CFG0                   ),
.RXDFE_GC_CFG1                   (RXDFE_GC_CFG1                   ),
.RXDFE_GC_CFG2                   (RXDFE_GC_CFG2                   ),
.RXDFE_H2_CFG0                   (RXDFE_H2_CFG0                   ),
.RXDFE_H2_CFG1                   (RXDFE_H2_CFG1                   ),
.RXDFE_H3_CFG0                   (RXDFE_H3_CFG0                   ),
.RXDFE_H3_CFG1                   (RXDFE_H3_CFG1                   ),
.RXDFE_H4_CFG0                   (RXDFE_H4_CFG0                   ),
.RXDFE_H4_CFG1                   (RXDFE_H4_CFG1                   ),
.RXDFE_H5_CFG0                   (RXDFE_H5_CFG0                   ),
.RXDFE_H5_CFG1                   (RXDFE_H5_CFG1                   ),
.RXDFE_H6_CFG0                   (RXDFE_H6_CFG0                   ),
.RXDFE_H6_CFG1                   (RXDFE_H6_CFG1                   ),
.RXDFE_H7_CFG0                   (RXDFE_H7_CFG0                   ),
.RXDFE_H7_CFG1                   (RXDFE_H7_CFG1                   ),
.RXDFE_H8_CFG0                   (RXDFE_H8_CFG0                   ),
.RXDFE_H8_CFG1                   (RXDFE_H8_CFG1                   ),
.RXDFE_H9_CFG0                   (RXDFE_H9_CFG0                   ),
.RXDFE_H9_CFG1                   (RXDFE_H9_CFG1                   ),
.RXDFE_HA_CFG0                   (RXDFE_HA_CFG0                   ),
.RXDFE_HA_CFG1                   (RXDFE_HA_CFG1                   ),
.RXDFE_HB_CFG0                   (RXDFE_HB_CFG0                   ),
.RXDFE_HB_CFG1                   (RXDFE_HB_CFG1                   ),
.RXDFE_HC_CFG0                   (RXDFE_HC_CFG0                   ),
.RXDFE_HC_CFG1                   (RXDFE_HC_CFG1                   ),
.RXDFE_HD_CFG0                   (RXDFE_HD_CFG0                   ),
.RXDFE_HD_CFG1                   (RXDFE_HD_CFG1                   ),
.RXDFE_HE_CFG0                   (RXDFE_HE_CFG0                   ),
.RXDFE_HE_CFG1                   (RXDFE_HE_CFG1                   ),
.RXDFE_HF_CFG0                   (RXDFE_HF_CFG0                   ),
.RXDFE_HF_CFG1                   (RXDFE_HF_CFG1                   ),
.RXDFE_KH_CFG0                   (RXDFE_KH_CFG0                   ),
.RXDFE_KH_CFG1                   (RXDFE_KH_CFG1                   ),
.RXDFE_KH_CFG2                   (RXDFE_KH_CFG2                   ),
.RXDFE_KH_CFG3                   (RXDFE_KH_CFG3                   ),
.RXDFE_OS_CFG0                   (RXDFE_OS_CFG0                   ),
.RXDFE_OS_CFG1                   (RXDFE_OS_CFG1                   ),
.RXDFE_UT_CFG0                   (RXDFE_UT_CFG0                   ),
.RXDFE_UT_CFG1                   (RXDFE_UT_CFG1                   ),
.RXDFE_UT_CFG2                   (RXDFE_UT_CFG2                   ),
.RXDFE_VP_CFG0                   (RXDFE_VP_CFG0                   ),
.RXDFE_VP_CFG1                   (RXDFE_VP_CFG1                   ),
.RXDLY_CFG                       (RXDLY_CFG                       ),
.RXDLY_LCFG                      (RXDLY_LCFG                      ),
.RXDLY_RAW_CFG                   (RXDLY_RAW_CFG                   ),
.RXDLY_RAW_LCFG                  (RXDLY_RAW_LCFG                  ),
.RXELECIDLE_CFG                  (RXELECIDLE_CFG                  ),
.RXGBOX_FIFO_INIT_RD_ADDR        (RXGBOX_FIFO_INIT_RD_ADDR        ),
.RXGEARBOX_EN                    (RXGEARBOX_EN                    ),
.RXISCANRESET_TIME               (RXISCANRESET_TIME               ),
.RXLPM_CFG                       (RXLPM_CFG                       ),
.RXLPM_GC_CFG                    (RXLPM_GC_CFG                    ),
.RXLPM_KH_CFG0                   (RXLPM_KH_CFG0                   ),
.RXLPM_KH_CFG1                   (RXLPM_KH_CFG1                   ),
.RXLPM_OS_CFG0                   (RXLPM_OS_CFG0                   ),
.RXLPM_OS_CFG1                   (RXLPM_OS_CFG1                   ),
.RXOSCALRESET_TIME               (RXOSCALRESET_TIME               ),
.RXOUT_DIV                       (RXOUT_DIV                       ),
.RXPCSRESET_TIME                 (RXPCSRESET_TIME                 ),
.RXPHBEACON_CFG                  (RXPHBEACON_CFG                  ),
.RXPHBEACON_RAW_CFG              (RXPHBEACON_RAW_CFG              ),
.RXPHDLY_CFG                     (RXPHDLY_CFG                     ),
.RXPHSAMP_CFG                    (RXPHSAMP_CFG                    ),
.RXPHSAMP_RAW_CFG                (RXPHSAMP_RAW_CFG                ),
.RXPHSLIP_CFG                    (RXPHSLIP_CFG                    ),
.RXPHSLIP_RAW_CFG                (RXPHSLIP_RAW_CFG                ),
.RXPH_MONITOR_SEL                (RXPH_MONITOR_SEL                ),
.RXPI_CFG0                       (RXPI_CFG0                       ),
.RXPI_CFG1                       (RXPI_CFG1                       ),
.RXPMACLK_SEL                    (RXPMACLK_SEL                    ),
.RXPMARESET_TIME                 (RXPMARESET_TIME                 ),
.RXPRBS_ERR_LOOPBACK             (RXPRBS_ERR_LOOPBACK             ),
.RXPRBS_LINKACQ_CNT              (RXPRBS_LINKACQ_CNT              ),
.RXRECCLKOUT0_SEL                (RXRECCLKOUT0_SEL                ),
.RXRECCLKOUT1_SEL                (RXRECCLKOUT1_SEL                ),
.RXREFCLKDIV2_SEL                (RXREFCLKDIV2_SEL                ),
.RXSLIDE_AUTO_WAIT               (RXSLIDE_AUTO_WAIT               ),
.RXSLIDE_MODE                    (RXSLIDE_MODE                    ),
.RXSYNC_MULTILANE                (RXSYNC_MULTILANE                ),
.RXSYNC_OVRD                     (RXSYNC_OVRD                     ),
.RXSYNC_SKIP_DA                  (RXSYNC_SKIP_DA                  ),
.RX_AFE_CM_EN                    (RX_AFE_CM_EN                    ),
.RX_BIAS_CFG0                    (RX_BIAS_CFG0                    ),
.RX_CAPFF_SARC_ENB               (RX_CAPFF_SARC_ENB               ),
.RX_CLK25_DIV                    (RX_CLK25_DIV                    ),
.RX_CLKMUX_EN                    (RX_CLKMUX_EN                    ),
.RX_CLK_SLIP_OVRD                (RX_CLK_SLIP_OVRD                ),
.RX_CM_BUF_CFG                   (RX_CM_BUF_CFG                   ),
.RX_CM_BUF_PD                    (RX_CM_BUF_PD                    ),
.RX_CM_SEL                       (RX_CM_SEL                       ),
.RX_CM_TRIM                      (RX_CM_TRIM                      ),
.RX_CTLE_PWR_SAVING              (RX_CTLE_PWR_SAVING              ),
.RX_CTLE_RES_CTRL                (RX_CTLE_RES_CTRL                ),
.RX_DATA_WIDTH                   (RX_DATA_WIDTH                   ),
.RX_DDI_SEL                      (RX_DDI_SEL                      ),
.RX_DEGEN_CTRL                   (RX_DEGEN_CTRL                   ),
.RX_DFELPM_CFG0                  (RX_DFELPM_CFG0                  ),
.RX_DFELPM_CFG1                  (RX_DFELPM_CFG1                  ),
.RX_DFELPM_KLKH_AGC_STUP_EN      (RX_DFELPM_KLKH_AGC_STUP_EN      ),
.RX_DFE_AGC_CFG1                 (RX_DFE_AGC_CFG1                 ),
.RX_DFE_KL_LPM_KH_CFG0           (RX_DFE_KL_LPM_KH_CFG0           ),
.RX_DFE_KL_LPM_KH_CFG1           (RX_DFE_KL_LPM_KH_CFG1           ),
.RX_DFE_KL_LPM_KL_CFG0           (RX_DFE_KL_LPM_KL_CFG0           ),
.RX_DFE_KL_LPM_KL_CFG1           (RX_DFE_KL_LPM_KL_CFG1           ),
.RX_DFE_LPM_HOLD_DURING_EIDLE    (RX_DFE_LPM_HOLD_DURING_EIDLE    ),
.RX_DISPERR_SEQ_MATCH            (RX_DISPERR_SEQ_MATCH            ),
.RX_DIVRESET_TIME                (RX_DIVRESET_TIME                ),
.RX_EN_CTLE_RCAL_B               (RX_EN_CTLE_RCAL_B               ),
.RX_EN_SUM_RCAL_B                (RX_EN_SUM_RCAL_B                ),
.RX_EYESCAN_VS_CODE              (RX_EYESCAN_VS_CODE              ),
.RX_EYESCAN_VS_NEG_DIR           (RX_EYESCAN_VS_NEG_DIR           ),
.RX_EYESCAN_VS_RANGE             (RX_EYESCAN_VS_RANGE             ),
.RX_EYESCAN_VS_UT_SIGN           (RX_EYESCAN_VS_UT_SIGN           ),
.RX_I2V_FILTER_EN                (RX_I2V_FILTER_EN                ),
.RX_INT_DATAWIDTH                (RX_INT_DATAWIDTH                ),
.RX_PMA_POWER_SAVE               (RX_PMA_POWER_SAVE               ),
.RX_PMA_RSV0                     (RX_PMA_RSV0                     ),
.RX_PROGDIV_CFG                  (RX_PROGDIV_CFG                  ),
.RX_PROGDIV_RATE                 (RX_PROGDIV_RATE                 ),
.RX_RESLOAD_CTRL                 (RX_RESLOAD_CTRL                 ),
.RX_RESLOAD_OVRD                 (RX_RESLOAD_OVRD                 ),
.RX_SAMPLE_PERIOD                (RX_SAMPLE_PERIOD                ),
.RX_SIG_VALID_DLY                (RX_SIG_VALID_DLY                ),
.RX_SUM_DEGEN_AVTT_OVERITE       (RX_SUM_DEGEN_AVTT_OVERITE       ),
.RX_SUM_DFETAPREP_EN             (RX_SUM_DFETAPREP_EN             ),
.RX_SUM_IREF_TUNE                (RX_SUM_IREF_TUNE                ),
.RX_SUM_PWR_SAVING               (RX_SUM_PWR_SAVING               ),
.RX_SUM_RES_CTRL                 (RX_SUM_RES_CTRL                 ),
.RX_SUM_VCMTUNE                  (RX_SUM_VCMTUNE                  ),
.RX_SUM_VCM_BIAS_TUNE_EN         (RX_SUM_VCM_BIAS_TUNE_EN         ),
.RX_SUM_VCM_OVWR                 (RX_SUM_VCM_OVWR                 ),
.RX_SUM_VREF_TUNE                (RX_SUM_VREF_TUNE                ),
.RX_TUNE_AFE_OS                  (RX_TUNE_AFE_OS                  ),
.RX_VREG_CTRL                    (RX_VREG_CTRL                    ),
.RX_VREG_PDB                     (RX_VREG_PDB                     ),
.RX_WIDEMODE_CDR                 (RX_WIDEMODE_CDR                 ),
.RX_WIDEMODE_CDR_GEN3            (RX_WIDEMODE_CDR_GEN3            ),
.RX_WIDEMODE_CDR_GEN4            (RX_WIDEMODE_CDR_GEN4            ),
.RX_XCLK_SEL                     (RX_XCLK_SEL                     ),
.RX_XMODE_SEL                    (RX_XMODE_SEL                    ),
.SAMPLE_CLK_PHASE                (SAMPLE_CLK_PHASE                ),
.SARC_ENB                        (SARC_ENB                        ),
.SARC_SEL                        (SARC_SEL                        ),
.SATA_CPLL_CFG                   (SATA_CPLL_CFG                   ),
.SDM0INITSEED0_0                 (SDM0INITSEED0_0                 ),
.SDM0INITSEED0_1                 (SDM0INITSEED0_1                 ),
.SDM1INITSEED0_0                 (SDM1INITSEED0_0                 ),
.SDM1INITSEED0_1                 (SDM1INITSEED0_1                 ),
.SIM_MODE                        (SIM_MODE                        ),
.SIM_RESET_SPEEDUP               (SIM_RESET_SPEEDUP               ),
.SIM_TX_EIDLE_DRIVE_LEVEL        (SIM_TX_EIDLE_DRIVE_LEVEL        ),
.SRSTMODE                        (SRSTMODE                        ),
.TAPDLY_SET_TX                   (TAPDLY_SET_TX                   ),
.TCO_NEW_CFG0                    (TCO_NEW_CFG0                    ),
.TCO_NEW_CFG1                    (TCO_NEW_CFG1                    ),
.TCO_NEW_CFG2                    (TCO_NEW_CFG2                    ),
.TCO_NEW_CFG3                    (TCO_NEW_CFG3                    ),
.TCO_RSVD1                       (TCO_RSVD1                       ),
.TCO_RSVD2                       (TCO_RSVD2                       ),
.TERM_RCAL_CFG                   (TERM_RCAL_CFG                   ),
.TERM_RCAL_OVRD                  (TERM_RCAL_OVRD                  ),
.TRANS_TIME_RATE                 (TRANS_TIME_RATE                 ),
.TST_RSV0                        (TST_RSV0                        ),
.TST_RSV1                        (TST_RSV1                        ),
.TXBUF_EN                        (TXBUF_EN                        ),
.TXDLY_CFG                       (TXDLY_CFG                       ),
.TXDLY_LCFG                      (TXDLY_LCFG                      ),
.TXDRV_FREQBAND                  (TXDRV_FREQBAND                  ),
.TXFE_CFG0                       (TXFE_CFG0                       ),
.TXFE_CFG1                       (TXFE_CFG1                       ),
.TXFE_CFG2                       (TXFE_CFG2                       ),
.TXFE_CFG3                       (TXFE_CFG3                       ),
.TXFIFO_ADDR_CFG                 (TXFIFO_ADDR_CFG                 ),
.TXGBOX_FIFO_INIT_RD_ADDR        (TXGBOX_FIFO_INIT_RD_ADDR        ),
.TXOUT_DIV                       (TXOUT_DIV                       ),
.TXPCSRESET_TIME                 (TXPCSRESET_TIME                 ),
.TXPHDLY_CFG0                    (TXPHDLY_CFG0                    ),
.TXPHDLY_CFG1                    (TXPHDLY_CFG1                    ),
.TXPH_CFG                        (TXPH_CFG                        ),
.TXPH_CFG2                       (TXPH_CFG2                       ),
.TXPH_MONITOR_SEL                (TXPH_MONITOR_SEL                ),
.TXPI_CFG0                       (TXPI_CFG0                       ),
.TXPI_CFG1                       (TXPI_CFG1                       ),
.TXPI_GRAY_SEL                   (TXPI_GRAY_SEL                   ),
.TXPI_INVSTROBE_SEL              (TXPI_INVSTROBE_SEL              ),
.TXPI_PPM                        (TXPI_PPM                        ),
.TXPI_PPM_CFG                    (TXPI_PPM_CFG                    ),
.TXPI_SYNFREQ_PPM                (TXPI_SYNFREQ_PPM                ),
.TXPMARESET_TIME                 (TXPMARESET_TIME                 ),
.TXREFCLKDIV2_SEL                (TXREFCLKDIV2_SEL                ),
.TXSWBST_BST                     (TXSWBST_BST                     ),
.TXSWBST_EN                      (TXSWBST_EN                      ),
.TXSWBST_MAG                     (TXSWBST_MAG                     ),
.TXSYNC_MULTILANE                (TXSYNC_MULTILANE                ),
.TXSYNC_OVRD                     (TXSYNC_OVRD                     ),
.TXSYNC_SKIP_DA                  (TXSYNC_SKIP_DA                  ),
.TX_CLK25_DIV                    (TX_CLK25_DIV                    ),
.TX_CLKMUX_EN                    (TX_CLKMUX_EN                    ),
.TX_DATA_WIDTH                   (TX_DATA_WIDTH                   ),
.TX_DCC_LOOP_RST_CFG             (TX_DCC_LOOP_RST_CFG             ),
.TX_DIVRESET_TIME                (TX_DIVRESET_TIME                ),
.TX_EIDLE_ASSERT_DELAY           (TX_EIDLE_ASSERT_DELAY           ),
.TX_EIDLE_DEASSERT_DELAY         (TX_EIDLE_DEASSERT_DELAY         ),
.TX_FABINT_USRCLK_FLOP           (TX_FABINT_USRCLK_FLOP           ),
.TX_FIFO_BYP_EN                  (TX_FIFO_BYP_EN                  ),
.TX_IDLE_DATA_ZERO               (TX_IDLE_DATA_ZERO               ),
.TX_INT_DATAWIDTH                (TX_INT_DATAWIDTH                ),
.TX_LOOPBACK_DRIVE_HIZ           (TX_LOOPBACK_DRIVE_HIZ           ),
.TX_MAINCURSOR_SEL               (TX_MAINCURSOR_SEL               ),
.TX_PHICAL_CFG0                  (TX_PHICAL_CFG0                  ),
.TX_PHICAL_CFG1                  (TX_PHICAL_CFG1                  ),
.TX_PI_BIASSET                   (TX_PI_BIASSET                   ),
.TX_PMADATA_OPT                  (TX_PMADATA_OPT                  ),
.TX_PMA_POWER_SAVE               (TX_PMA_POWER_SAVE               ),
.TX_PMA_RSV0                     (TX_PMA_RSV0                     ),
.TX_PMA_RSV1                     (TX_PMA_RSV1                     ),
.TX_PROGCLK_SEL                  (TX_PROGCLK_SEL                  ),
.TX_PROGDIV_CFG                  (TX_PROGDIV_CFG                  ),
.TX_PROGDIV_RATE                 (TX_PROGDIV_RATE                 ),
.TX_SAMPLE_PERIOD                (TX_SAMPLE_PERIOD                ),
.TX_SW_MEAS                      (TX_SW_MEAS                      ),
.TX_VREG_CTRL                    (TX_VREG_CTRL                    ),
.TX_VREG_PDB                     (TX_VREG_PDB                     ),
.TX_VREG_VREFSEL                 (TX_VREG_VREFSEL                 ),
.TX_XCLK_SEL                     (TX_XCLK_SEL                     ),
.USE_PCS_CLK_PHASE_SEL           (USE_PCS_CLK_PHASE_SEL           ),
.USE_RAW_ELEC                    (USE_RAW_ELEC                    ),
.Y_ALL_MODE                      (Y_ALL_MODE                      )
) inst (
.gtwiz_reset_clk_freerun_in           (gtwiz_reset_clk_freerun_in           ),
.gtwiz_reset_all_in                   (gtwiz_reset_all_in                   ),
.gtwiz_reset_tx_pll_and_datapath_in   (gtwiz_reset_tx_pll_and_datapath_in   ),
.gtwiz_reset_tx_datapath_in           (gtwiz_reset_tx_datapath_in           ),
.gtwiz_reset_rx_pll_and_datapath_in   (gtwiz_reset_rx_pll_and_datapath_in   ),
.gtwiz_reset_rx_datapath_in           (gtwiz_reset_rx_datapath_in           ),
.gtwiz_reset_rx_cdr_stable_out        (gtwiz_reset_rx_cdr_stable_out        ),
.gtwiz_reset_tx_done_out              (gtwiz_reset_tx_done_out              ),
.gtwiz_reset_rx_done_out              (gtwiz_reset_rx_done_out              ),
.gtwiz_pllreset_rx_out                (gtwiz_pllreset_rx_out                ),
.gtwiz_pllreset_tx_out                (gtwiz_pllreset_tx_out                ),
.plllock_tx_in                        (plllock_tx_in                        ),
.plllock_rx_in                        (plllock_rx_in                        ),
.gtf_ch_cdrstepdir                    (gtf_ch_cdrstepdir                    ),
.gtf_ch_cdrstepsq                     (gtf_ch_cdrstepsq                     ),
.gtf_ch_cdrstepsx                     (gtf_ch_cdrstepsx                     ),
.gtf_ch_cfgreset                      (gtf_ch_cfgreset                      ),
.gtf_ch_clkrsvd0                      (gtf_ch_clkrsvd0                      ),
.gtf_ch_clkrsvd1                      (gtf_ch_clkrsvd1                      ),
.gtf_ch_cpllfreqlock                  (gtf_ch_cpllfreqlock                  ),
.gtf_ch_cplllockdetclk                (gtf_ch_cplllockdetclk                ),
.gtf_ch_cplllocken                    (gtf_ch_cplllocken                    ),
.gtf_ch_cpllpd                        (gtf_ch_cpllpd                        ),
.gtf_ch_cpllreset                     (gtf_ch_cpllreset                     ),
.gtf_ch_ctltxresendpause              (gtf_ch_ctltxresendpause              ),
.gtf_ch_dmonfiforeset                 (gtf_ch_dmonfiforeset                 ),
.gtf_ch_dmonitorclk                   (gtf_ch_dmonitorclk                   ),
.gtf_ch_drpclk                        (gtf_ch_drpclk                        ),
.gtf_ch_drprst                        (gtf_ch_drprst                        ),
.gtf_ch_eyescanreset                  (gtf_ch_eyescanreset                  ),
.gtf_ch_eyescantrigger                (gtf_ch_eyescantrigger                ),
.gtf_ch_freqos                        (gtf_ch_freqos                        ),
.gtf_ch_gtfrxn                        (gtf_ch_gtfrxn                        ),
.gtf_ch_gtfrxp                        (gtf_ch_gtfrxp                        ),
.gtf_ch_gtgrefclk                     (gtf_ch_gtgrefclk                     ),
.gtf_ch_gtnorthrefclk0                (gtf_ch_gtnorthrefclk0                ),
.gtf_ch_gtnorthrefclk1                (gtf_ch_gtnorthrefclk1                ),
.gtf_ch_gtrefclk0                     (gtf_ch_gtrefclk0                     ),
.gtf_ch_gtrefclk1                     (gtf_ch_gtrefclk1                     ),
.gtf_ch_gtrxresetsel                  (gtf_ch_gtrxresetsel                  ),
.gtf_ch_gtsouthrefclk0                (gtf_ch_gtsouthrefclk0                ),
.gtf_ch_gtsouthrefclk1                (gtf_ch_gtsouthrefclk1                ),
.gtf_ch_gttxresetsel                  (gtf_ch_gttxresetsel                  ),
.gtf_ch_incpctrl                      (gtf_ch_incpctrl                      ),
.gtf_ch_qpll0clk                      (gtf_ch_qpll0clk                      ),
.gtf_ch_qpll0freqlock                 (gtf_ch_qpll0freqlock                 ),
.gtf_ch_qpll0refclk                   (gtf_ch_qpll0refclk                   ),
.gtf_ch_qpll1clk                      (gtf_ch_qpll1clk                      ),
.gtf_ch_qpll1freqlock                 (gtf_ch_qpll1freqlock                 ),
.gtf_ch_qpll1refclk                   (gtf_ch_qpll1refclk                   ),
.gtf_ch_resetovrd                     (gtf_ch_resetovrd                     ),
.gtf_ch_rxafecfoken                   (gtf_ch_rxafecfoken                   ),
.gtf_ch_rxcdrfreqreset                (gtf_ch_rxcdrfreqreset                ),
.gtf_ch_rxcdrhold                     (gtf_ch_rxcdrhold                     ),
.gtf_ch_rxcdrovrden                   (gtf_ch_rxcdrovrden                   ),
.gtf_ch_rxcdrreset                    (gtf_ch_rxcdrreset                    ),
.gtf_ch_rxckcalreset                  (gtf_ch_rxckcalreset                  ),
.gtf_ch_rxdfeagchold                  (gtf_ch_rxdfeagchold                  ),
.gtf_ch_rxdfeagcovrden                (gtf_ch_rxdfeagcovrden                ),
.gtf_ch_rxdfecfokfen                  (gtf_ch_rxdfecfokfen                  ),
.gtf_ch_rxdfecfokfpulse               (gtf_ch_rxdfecfokfpulse               ),
.gtf_ch_rxdfecfokhold                 (gtf_ch_rxdfecfokhold                 ),
.gtf_ch_rxdfecfokovren                (gtf_ch_rxdfecfokovren                ),
.gtf_ch_rxdfekhhold                   (gtf_ch_rxdfekhhold                   ),
.gtf_ch_rxdfekhovrden                 (gtf_ch_rxdfekhovrden                 ),
.gtf_ch_rxdfelfhold                   (gtf_ch_rxdfelfhold                   ),
.gtf_ch_rxdfelfovrden                 (gtf_ch_rxdfelfovrden                 ),
.gtf_ch_rxdfelpmreset                 (gtf_ch_rxdfelpmreset                 ),
.gtf_ch_rxdfetap10hold                (gtf_ch_rxdfetap10hold                ),
.gtf_ch_rxdfetap10ovrden              (gtf_ch_rxdfetap10ovrden              ),
.gtf_ch_rxdfetap11hold                (gtf_ch_rxdfetap11hold                ),
.gtf_ch_rxdfetap11ovrden              (gtf_ch_rxdfetap11ovrden              ),
.gtf_ch_rxdfetap12hold                (gtf_ch_rxdfetap12hold                ),
.gtf_ch_rxdfetap12ovrden              (gtf_ch_rxdfetap12ovrden              ),
.gtf_ch_rxdfetap13hold                (gtf_ch_rxdfetap13hold                ),
.gtf_ch_rxdfetap13ovrden              (gtf_ch_rxdfetap13ovrden              ),
.gtf_ch_rxdfetap14hold                (gtf_ch_rxdfetap14hold                ),
.gtf_ch_rxdfetap14ovrden              (gtf_ch_rxdfetap14ovrden              ),
.gtf_ch_rxdfetap15hold                (gtf_ch_rxdfetap15hold                ),
.gtf_ch_rxdfetap15ovrden              (gtf_ch_rxdfetap15ovrden              ),
.gtf_ch_rxdfetap2hold                 (gtf_ch_rxdfetap2hold                 ),
.gtf_ch_rxdfetap2ovrden               (gtf_ch_rxdfetap2ovrden               ),
.gtf_ch_rxdfetap3hold                 (gtf_ch_rxdfetap3hold                 ),
.gtf_ch_rxdfetap3ovrden               (gtf_ch_rxdfetap3ovrden               ),
.gtf_ch_rxdfetap4hold                 (gtf_ch_rxdfetap4hold                 ),
.gtf_ch_rxdfetap4ovrden               (gtf_ch_rxdfetap4ovrden               ),
.gtf_ch_rxdfetap5hold                 (gtf_ch_rxdfetap5hold                 ),
.gtf_ch_rxdfetap5ovrden               (gtf_ch_rxdfetap5ovrden               ),
.gtf_ch_rxdfetap6hold                 (gtf_ch_rxdfetap6hold                 ),
.gtf_ch_rxdfetap6ovrden               (gtf_ch_rxdfetap6ovrden               ),
.gtf_ch_rxdfetap7hold                 (gtf_ch_rxdfetap7hold                 ),
.gtf_ch_rxdfetap7ovrden               (gtf_ch_rxdfetap7ovrden               ),
.gtf_ch_rxdfetap8hold                 (gtf_ch_rxdfetap8hold                 ),
.gtf_ch_rxdfetap8ovrden               (gtf_ch_rxdfetap8ovrden               ),
.gtf_ch_rxdfetap9hold                 (gtf_ch_rxdfetap9hold                 ),
.gtf_ch_rxdfetap9ovrden               (gtf_ch_rxdfetap9ovrden               ),
.gtf_ch_rxdfeuthold                   (gtf_ch_rxdfeuthold                   ),
.gtf_ch_rxdfeutovrden                 (gtf_ch_rxdfeutovrden                 ),
.gtf_ch_rxdfevphold                   (gtf_ch_rxdfevphold                   ),
.gtf_ch_rxdfevpovrden                 (gtf_ch_rxdfevpovrden                 ),
.gtf_ch_rxdfexyden                    (gtf_ch_rxdfexyden                    ),




.gtf_ch_rxlpmen                       (gtf_ch_rxlpmen                       ),
.gtf_ch_rxlpmgchold                   (gtf_ch_rxlpmgchold                   ),
.gtf_ch_rxlpmgcovrden                 (gtf_ch_rxlpmgcovrden                 ),
.gtf_ch_rxlpmhfhold                   (gtf_ch_rxlpmhfhold                   ),
.gtf_ch_rxlpmhfovrden                 (gtf_ch_rxlpmhfovrden                 ),
.gtf_ch_rxlpmlfhold                   (gtf_ch_rxlpmlfhold                   ),
.gtf_ch_rxlpmlfklovrden               (gtf_ch_rxlpmlfklovrden               ),
.gtf_ch_rxlpmoshold                   (gtf_ch_rxlpmoshold                   ),
.gtf_ch_rxlpmosovrden                 (gtf_ch_rxlpmosovrden                 ),
.gtf_ch_rxoscalreset                  (gtf_ch_rxoscalreset                  ),
.gtf_ch_rxoshold                      (gtf_ch_rxoshold                      ),
.gtf_ch_rxosovrden                    (gtf_ch_rxosovrden                    ),
.gtf_ch_rxpcsreset                    (gtf_ch_rxpcsreset                    ),
.gtf_ch_rxslippma                     (gtf_ch_rxslippma                     ),



.gtwiz_buffbypass_rx_done_out         (gtwiz_buffbypass_rx_done_out         ),
.gtf_ch_rxpmareset                    (gtf_ch_rxpmareset                    ),
.gtf_ch_rxpolarity                    (gtf_ch_rxpolarity                    ),
.gtf_ch_rxprbscntreset                (gtf_ch_rxprbscntreset                ),
.gtf_ch_rxslipoutclk                  (gtf_ch_rxslipoutclk                  ),



.gtf_ch_rxtermination                 (gtf_ch_rxtermination                 ),
.gtf_ch_rxuserrdy                     (gtf_ch_rxuserrdy                     ),
.gtf_ch_txaxisterr                    (gtf_ch_txaxisterr                    ),
.gtf_ch_txaxistpoison                 (gtf_ch_txaxistpoison                 ),
.gtf_ch_txaxistvalid                  (gtf_ch_txaxistvalid                  ),
.gtf_ch_txdccforcestart               (gtf_ch_txdccforcestart               ),
.gtf_ch_txdccreset                    (gtf_ch_txdccreset                    ),
.gtf_ch_txelecidle                    (gtf_ch_txelecidle                    ),
.gtf_ch_txgbseqsync                   (gtf_ch_txgbseqsync                   ),
.gtf_ch_txmuxdcdexhold                (gtf_ch_txmuxdcdexhold                ),
.gtf_ch_txmuxdcdorwren                (gtf_ch_txmuxdcdorwren                ),
.gtf_ch_txpcsreset                    (gtf_ch_txpcsreset                    ),
.gtf_ch_txpippmen                     (gtf_ch_txpippmen                     ),
.gtf_ch_txpippmovrden                 (gtf_ch_txpippmovrden                 ),
.gtf_ch_txpippmpd                     (gtf_ch_txpippmpd                     ),
.gtf_ch_txpippmsel                    (gtf_ch_txpippmsel                    ),
.gtf_ch_txpisopd                      (gtf_ch_txpisopd                      ),
.gtf_ch_txpmareset                    (gtf_ch_txpmareset                    ),
.gtf_ch_txpolarity                    (gtf_ch_txpolarity                    ),
.gtf_ch_txprbsforceerr                (gtf_ch_txprbsforceerr                ),
.gtf_ch_txuserrdy                     (gtf_ch_txuserrdy                     ),
.gtf_ch_gtrsvd                        (gtf_ch_gtrsvd                        ),
.gtf_ch_pcsrsvdin                     (gtf_ch_pcsrsvdin                     ),
.gtf_ch_tstin                         (gtf_ch_tstin                         ),
.gtf_ch_rxelecidlemode                (gtf_ch_rxelecidlemode                ),
.gtf_ch_rxmonitorsel                  (gtf_ch_rxmonitorsel                  ),
.gtf_ch_rxpd                          (gtf_ch_rxpd                          ),
.gtf_ch_rxpllclksel                   (gtf_ch_rxpllclksel                   ),
.gtf_ch_rxsysclksel                   (gtf_ch_rxsysclksel                   ),
.gtf_ch_txaxistsof                    (gtf_ch_txaxistsof                    ),
.gtf_ch_txpd                          (gtf_ch_txpd                          ),
.gtf_ch_txpllclksel                   (gtf_ch_txpllclksel                   ),
.gtf_ch_txsysclksel                   (gtf_ch_txsysclksel                   ),
.gtf_ch_cpllrefclksel                 (gtf_ch_cpllrefclksel                 ),
.gtf_ch_rxoutclksel                   (gtf_ch_rxoutclksel                   ),
.gtf_ch_txoutclksel                   (gtf_ch_txoutclksel                   ),
.gtf_ch_txrawdata                     (gtf_ch_txrawdata                     ),
.gtf_ch_rxdfecfokfcnum                (gtf_ch_rxdfecfokfcnum                ),
.gtf_ch_rxprbssel                     (gtf_ch_rxprbssel                     ),
.gtf_ch_txprbssel                     (gtf_ch_txprbssel                     ),
.gtf_ch_txaxistterm                   (gtf_ch_txaxistterm                   ),
.gtf_ch_txdiffctrl                    (gtf_ch_txdiffctrl                    ),
.gtf_ch_txpippmstepsize               (gtf_ch_txpippmstepsize               ),
.gtf_ch_txpostcursor                  (gtf_ch_txpostcursor                  ),
.gtf_ch_txprecursor                   (gtf_ch_txprecursor                   ),
.gtf_ch_txaxistdata                   (gtf_ch_txaxistdata                   ),
.gtf_ch_rxckcalstart                  (gtf_ch_rxckcalstart                  ),
.gtf_ch_txmaincursor                  (gtf_ch_txmaincursor                  ),
.gtf_ch_txaxistlast                   (gtf_ch_txaxistlast                   ),
.gtf_ch_txaxistpre                    (gtf_ch_txaxistpre                    ),
.gtf_ch_ctlrxpauseack                 (gtf_ch_ctlrxpauseack                 ),
.gtf_ch_ctltxpausereq                 (gtf_ch_ctltxpausereq                 ),
.gtf_ch_cpllfbclklost                 (gtf_ch_cpllfbclklost                 ),
.gtf_ch_cplllock                      (gtf_ch_cplllock                      ),
.gtf_ch_cpllrefclklost                (gtf_ch_cpllrefclklost                ),
.gtf_ch_dmonitoroutclk                (gtf_ch_dmonitoroutclk                ),
.gtf_ch_eyescandataerror              (gtf_ch_eyescandataerror              ),
.gtf_ch_gtftxn                        (gtf_ch_gtftxn                        ),
.gtf_ch_gtftxp                        (gtf_ch_gtftxp                        ),
.gtf_ch_gtpowergood                   (gtf_ch_gtpowergood                   ),
.gtf_ch_gtrefclkmonitor               (gtf_ch_gtrefclkmonitor               ),
.gtf_ch_resetexception                (gtf_ch_resetexception                ),
.gtf_ch_rxaxisterr                    (gtf_ch_rxaxisterr                    ),
.gtf_ch_rxaxistvalid                  (gtf_ch_rxaxistvalid                  ),
.gtf_ch_rxbitslip                     (gtf_ch_rxbitslip                     ),
.gtf_ch_rxcdrlock                     (gtf_ch_rxcdrlock                     ),
.gtf_ch_rxcdrphdone                   (gtf_ch_rxcdrphdone                   ),
.gtf_ch_rxckcaldone                   (gtf_ch_rxckcaldone                   ),

.gtf_ch_rxelecidle                    (gtf_ch_rxelecidle                    ),
.gtf_ch_rxgbseqstart                  (gtf_ch_rxgbseqstart                  ),
.gtf_ch_rxosintdone                   (gtf_ch_rxosintdone                   ),
.gtf_ch_rxosintstarted                (gtf_ch_rxosintstarted                ),
.gtf_ch_rxosintstrobedone             (gtf_ch_rxosintstrobedone             ),
.gtf_ch_rxosintstrobestarted          (gtf_ch_rxosintstrobestarted          ),
.gtf_ch_rxoutclk                      (gtf_ch_rxoutclk                      ),
.gtf_ch_rxoutclkfabric                (gtf_ch_rxoutclkfabric                ),
.gtf_ch_rxoutclkpcs                   (gtf_ch_rxoutclkpcs                   ),

.gtf_ch_rxphalignerr                  (gtf_ch_rxphalignerr                  ),
.gtf_ch_rxpmaresetdone                (gtf_ch_rxpmaresetdone                ),
.gtf_ch_rxprbserr                     (gtf_ch_rxprbserr                     ),
.gtf_ch_rxprbslocked                  (gtf_ch_rxprbslocked                  ),
.gtf_ch_rxprgdivresetdone             (gtf_ch_rxprgdivresetdone             ),
.gtf_ch_rxptpsop                      (gtf_ch_rxptpsop                      ),
.gtf_ch_rxptpsoppos                   (gtf_ch_rxptpsoppos                   ),
.gtf_ch_rxrecclkout                   (gtf_ch_rxrecclkout                   ),
.gtf_ch_rxresetdone                   (gtf_ch_rxresetdone                   ),
.gtf_ch_rxslipdone                    (gtf_ch_rxslipdone                    ),
.gtf_ch_rxslipoutclkrdy               (gtf_ch_rxslipoutclkrdy               ),
.gtf_ch_rxslippmardy                  (gtf_ch_rxslippmardy                  ),
.gtf_ch_rxsyncdone                    (gtf_ch_rxsyncdone                    ),





.gtf_ch_statrxblocklock               (gtf_ch_statrxblocklock               ),

.gtf_ch_statrxfcserr                  (gtf_ch_statrxfcserr                  ),

.gtf_ch_ctltxsendidle                 (gtf_ch_ctltxsendidle                 ),
.gtf_ch_ctltxsendlfi                  (gtf_ch_ctltxsendlfi                  ),
.gtf_ch_ctltxsendrfi                  (gtf_ch_ctltxsendrfi                  ),

.gtf_ch_loopback                      (gtf_ch_loopback                      ),
.gtf_ch_statrxhiber                   (gtf_ch_statrxhiber                   ),
.gtf_ch_statrxstatus                  (gtf_ch_statrxstatus                  ),
.gtf_ch_statrxpkterr                  (gtf_ch_statrxpkterr                  ),
.gtf_ch_statrxbadpreamble             (gtf_ch_statrxbadpreamble             ),
.gtf_ch_statrxbadsfd                  (gtf_ch_statrxbadsfd                  ),
.gtf_ch_statrxgotsignalos             (gtf_ch_statrxgotsignalos             ),
.gtf_ch_statrxbadcode                 (gtf_ch_statrxbadcode                 ),
.gtf_ch_statrxstompedfcs              (gtf_ch_statrxstompedfcs              ),
.gtf_ch_statrxframingerr              (gtf_ch_statrxframingerr              ),
.gtf_ch_statrxtruncated               (gtf_ch_statrxtruncated               ),
.gtf_ch_statrxbytes                   (gtf_ch_statrxbytes                   ),
.gtf_ch_statrxpkt                     (gtf_ch_statrxpkt                     ),
.gtf_ch_statrxbadfcs                  (gtf_ch_statrxbadfcs                  ),
.gtf_ch_statrxunicast                 (gtf_ch_statrxunicast                 ),
.gtf_ch_statrxbroadcast               (gtf_ch_statrxbroadcast               ),
.gtf_ch_statrxvlan                    (gtf_ch_statrxvlan                    ),
.gtf_ch_statrxinrangeerr              (gtf_ch_statrxinrangeerr              ),
.gtf_ch_statrxpausevalid              (gtf_ch_statrxpausevalid              ),
.gtf_ch_statrxpausereq                (gtf_ch_statrxpausereq                ),
.gtf_ch_statrxpausequanta             (gtf_ch_statrxpausequanta             ),
.gtf_ch_stattxbytes                   (gtf_ch_stattxbytes                   ),
.gtf_ch_stattxpkt                     (gtf_ch_stattxpkt                     ),
.gtf_ch_stattxpkterr                  (gtf_ch_stattxpkterr                  ),
.gtf_ch_stattxbadfcs                  (gtf_ch_stattxbadfcs                  ),
.gtf_ch_stattxunicast                 (gtf_ch_stattxunicast                 ),
.gtf_ch_stattxbroadcast               (gtf_ch_stattxbroadcast               ),
.gtf_ch_stattxmulticast               (gtf_ch_stattxmulticast               ),
.gtf_ch_stattxvlan                    (gtf_ch_stattxvlan                    ),
.gtf_ch_statrxmulticast               (gtf_ch_statrxmulticast               ),
.gtf_ch_statrxinternallocalfault      (gtf_ch_statrxinternallocalfault      ),
.gtf_ch_statrxlocalfault              (gtf_ch_statrxlocalfault              ),
.gtf_ch_statrxreceivedlocalfault      (gtf_ch_statrxreceivedlocalfault      ),
.gtf_ch_statrxremotefault             (gtf_ch_statrxremotefault             ),
.gtf_ch_statrxtestpatternmismatch     (gtf_ch_statrxtestpatternmismatch     ),
.gtf_ch_statrxvalidctrlcode           (gtf_ch_statrxvalidctrlcode           ),
.gtf_ch_stattxfcserr                  (gtf_ch_stattxfcserr                  ),
.gtf_ch_txaxistready                  (gtf_ch_txaxistready                  ),
.gtf_ch_txdccdone                     (gtf_ch_txdccdone                     ),
.gtf_ch_txgbseqstart                  (gtf_ch_txgbseqstart                  ),
.gtf_ch_txoutclk                      (gtf_ch_txoutclk                      ),
.gtf_ch_txoutclkfabric                (gtf_ch_txoutclkfabric                ),
.gtf_ch_txoutclkpcs                   (gtf_ch_txoutclkpcs                   ),
.gtf_ch_txpmaresetdone                (gtf_ch_txpmaresetdone                ),
.gtf_ch_txprgdivresetdone             (gtf_ch_txprgdivresetdone             ),
.gtf_ch_txptpsop                      (gtf_ch_txptpsop                      ),
.gtf_ch_txptpsoppos                   (gtf_ch_txptpsoppos                   ),
.gtf_ch_txresetdone                   (gtf_ch_txresetdone                   ),
.gtf_ch_txsyncdone                    (gtf_ch_txsyncdone                    ),
.gtf_ch_txunfout                      (gtf_ch_txunfout                      ),
.gtf_ch_txaxistcanstart               (gtf_ch_txaxistcanstart               ),
.gtf_ch_rxinvalidstart                (gtf_ch_rxinvalidstart                ),
.gtf_ch_pcsrsvdout                    (gtf_ch_pcsrsvdout                    ),
.gtf_ch_pinrsrvdas                    (gtf_ch_pinrsrvdas                    ),
.gtf_ch_rxaxistsof                    (gtf_ch_rxaxistsof                    ),
.gtf_ch_rxrawdata                     (gtf_ch_rxrawdata                     ),


.gtf_ch_rxaxistterm                   (gtf_ch_rxaxistterm                   ),
.gtf_ch_rxaxistdata                   (gtf_ch_rxaxistdata                   ),
.gtf_ch_rxaxistlast                   (gtf_ch_rxaxistlast                   ),
.gtf_ch_rxaxistpre                    (gtf_ch_rxaxistpre                    ),
.gtf_ch_rxmonitorout                  (gtf_ch_rxmonitorout                  ),



.gtf_ch_stattxpausevalid              (gtf_ch_stattxpausevalid              ),
.gtf_ch_gttxreset_out                 (gtf_ch_gttxreset_out                 ),
 .gtwiz_buffbypass_tx_done_out        (gtwiz_buffbypass_tx_done_out         ),
.gtf_txusrclk2_out                    (gtf_txusrclk2_out                    ),
.gtf_rxusrclk2_out                    (gtf_rxusrclk2_out                    )
);
endmodule
`default_nettype wire
//------}
